VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO address_gen
  CLASS BLOCK ;
  FOREIGN address_gen ;
  ORIGIN 1.900 4.000 ;
  SIZE 199.000 BY 188.300 ;
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 1.200 161.600 2.000 170.200 ;
        RECT 4.400 161.600 5.200 170.200 ;
        RECT 7.600 161.600 8.400 170.200 ;
        RECT 10.800 161.600 11.600 170.200 ;
        RECT 14.000 161.600 14.800 170.200 ;
        RECT 17.200 161.600 18.000 170.200 ;
        RECT 22.800 161.600 23.600 166.200 ;
        RECT 26.000 161.600 26.800 166.200 ;
        RECT 31.600 161.600 32.400 170.000 ;
        RECT 36.400 161.600 37.200 169.000 ;
        RECT 41.200 161.600 42.000 170.000 ;
        RECT 46.800 161.600 47.600 166.200 ;
        RECT 50.000 161.600 50.800 166.200 ;
        RECT 55.600 161.600 56.400 170.200 ;
        RECT 65.200 161.600 66.000 169.000 ;
        RECT 70.000 161.600 70.800 169.000 ;
        RECT 74.800 161.600 75.600 169.000 ;
        RECT 79.600 161.600 80.400 170.200 ;
        RECT 85.200 161.600 86.000 166.200 ;
        RECT 88.400 161.600 89.200 166.200 ;
        RECT 94.000 161.600 94.800 170.000 ;
        RECT 98.800 161.600 99.600 169.000 ;
        RECT 103.600 161.600 104.400 169.000 ;
        RECT 108.400 161.600 109.200 170.200 ;
        RECT 114.000 161.600 114.800 166.200 ;
        RECT 117.200 161.600 118.000 166.200 ;
        RECT 122.800 161.600 123.600 170.000 ;
        RECT 127.600 161.600 128.400 169.000 ;
        RECT 132.400 161.600 133.200 169.000 ;
        RECT 142.000 161.600 142.800 170.200 ;
        RECT 147.600 161.600 148.400 166.200 ;
        RECT 150.800 161.600 151.600 166.200 ;
        RECT 156.400 161.600 157.200 170.000 ;
        RECT 161.200 161.600 162.000 169.000 ;
        RECT 166.000 161.600 166.800 170.000 ;
        RECT 171.600 161.600 172.400 166.200 ;
        RECT 174.800 161.600 175.600 166.200 ;
        RECT 180.400 161.600 181.200 170.200 ;
        RECT 185.800 161.600 186.600 170.200 ;
        RECT 191.600 161.600 192.400 169.000 ;
        RECT 0.400 160.400 194.800 161.600 ;
        RECT 2.800 151.800 3.600 160.400 ;
        RECT 8.400 155.800 9.200 160.400 ;
        RECT 11.600 155.800 12.400 160.400 ;
        RECT 17.200 152.000 18.000 160.400 ;
        RECT 22.000 151.800 22.800 160.400 ;
        RECT 27.600 155.800 28.400 160.400 ;
        RECT 30.800 155.800 31.600 160.400 ;
        RECT 36.400 152.000 37.200 160.400 ;
        RECT 41.200 152.200 42.000 160.400 ;
        RECT 44.400 155.800 45.200 160.400 ;
        RECT 46.000 155.800 46.800 160.400 ;
        RECT 50.800 153.000 51.600 160.400 ;
        RECT 60.400 155.800 61.200 160.400 ;
        RECT 63.600 155.800 64.400 160.400 ;
        RECT 65.200 155.800 66.000 160.400 ;
        RECT 71.600 153.000 72.400 160.400 ;
        RECT 74.800 155.800 75.600 160.400 ;
        RECT 78.000 155.800 78.800 160.400 ;
        RECT 79.600 155.800 80.400 160.400 ;
        RECT 85.000 151.800 85.800 160.400 ;
        RECT 90.800 153.000 91.600 160.400 ;
        RECT 95.600 155.800 96.400 160.400 ;
        RECT 98.800 152.200 99.600 160.400 ;
        RECT 102.000 151.800 102.800 160.400 ;
        RECT 105.200 151.800 106.000 160.400 ;
        RECT 108.400 151.800 109.200 160.400 ;
        RECT 111.600 151.800 112.400 160.400 ;
        RECT 114.800 151.800 115.600 160.400 ;
        RECT 118.000 153.000 118.800 160.400 ;
        RECT 123.400 155.800 124.200 160.400 ;
        RECT 127.600 151.800 128.400 160.400 ;
        RECT 129.200 155.800 130.000 160.400 ;
        RECT 132.400 155.800 133.200 160.400 ;
        RECT 140.400 153.000 141.200 160.400 ;
        RECT 145.200 151.800 146.000 160.400 ;
        RECT 149.400 155.800 150.200 160.400 ;
        RECT 154.800 151.800 155.600 160.400 ;
        RECT 158.000 151.800 158.800 160.400 ;
        RECT 163.600 155.800 164.400 160.400 ;
        RECT 166.800 155.800 167.600 160.400 ;
        RECT 172.400 152.000 173.200 160.400 ;
        RECT 177.200 152.000 178.000 160.400 ;
        RECT 182.800 155.800 183.600 160.400 ;
        RECT 186.000 155.800 186.800 160.400 ;
        RECT 191.600 151.800 192.400 160.400 ;
        RECT 2.800 121.600 3.600 129.000 ;
        RECT 7.600 121.600 8.400 129.000 ;
        RECT 12.400 121.600 13.200 129.000 ;
        RECT 17.200 121.600 18.000 130.200 ;
        RECT 21.400 121.600 22.200 126.200 ;
        RECT 23.600 121.600 24.400 126.200 ;
        RECT 26.800 121.600 27.600 126.200 ;
        RECT 30.000 121.600 30.800 126.200 ;
        RECT 33.800 121.600 34.600 130.200 ;
        RECT 39.600 121.600 40.400 129.000 ;
        RECT 47.600 121.600 48.400 130.200 ;
        RECT 50.800 121.600 51.600 126.200 ;
        RECT 58.800 121.600 59.600 129.000 ;
        RECT 63.600 121.600 64.400 126.200 ;
        RECT 66.800 121.600 67.600 126.200 ;
        RECT 69.000 121.600 69.800 126.200 ;
        RECT 73.200 121.600 74.000 130.200 ;
        RECT 78.000 121.600 78.800 130.200 ;
        RECT 79.600 121.600 80.400 126.200 ;
        RECT 82.800 121.600 83.600 126.200 ;
        RECT 86.000 121.600 86.800 130.200 ;
        RECT 91.600 121.600 92.400 126.200 ;
        RECT 94.800 121.600 95.600 126.200 ;
        RECT 100.400 121.600 101.200 130.000 ;
        RECT 105.200 121.600 106.000 130.200 ;
        RECT 110.800 121.600 111.600 126.200 ;
        RECT 114.000 121.600 114.800 126.200 ;
        RECT 119.600 121.600 120.400 130.000 ;
        RECT 122.800 121.600 123.600 130.200 ;
        RECT 127.600 121.600 128.400 126.200 ;
        RECT 130.800 121.600 131.600 126.200 ;
        RECT 135.600 121.600 136.400 129.000 ;
        RECT 143.600 121.600 144.400 126.200 ;
        RECT 146.800 121.600 147.600 130.200 ;
        RECT 153.200 121.600 154.000 129.000 ;
        RECT 158.000 121.600 158.800 130.200 ;
        RECT 162.200 121.600 163.000 126.200 ;
        RECT 164.400 121.600 165.200 126.200 ;
        RECT 167.600 121.600 168.400 126.200 ;
        RECT 172.400 121.600 173.200 129.000 ;
        RECT 177.200 121.600 178.000 130.000 ;
        RECT 182.800 121.600 183.600 126.200 ;
        RECT 186.000 121.600 186.800 126.200 ;
        RECT 191.600 121.600 192.400 130.200 ;
        RECT 0.400 120.400 194.800 121.600 ;
        RECT 2.800 113.000 3.600 120.400 ;
        RECT 7.600 111.800 8.400 120.400 ;
        RECT 13.200 115.800 14.000 120.400 ;
        RECT 16.400 115.800 17.200 120.400 ;
        RECT 22.000 112.000 22.800 120.400 ;
        RECT 26.800 112.200 27.600 120.400 ;
        RECT 30.000 115.800 30.800 120.400 ;
        RECT 31.600 115.800 32.400 120.400 ;
        RECT 34.800 111.800 35.600 120.400 ;
        RECT 39.600 111.800 40.400 120.400 ;
        RECT 43.800 115.800 44.600 120.400 ;
        RECT 47.600 116.200 48.400 120.400 ;
        RECT 50.800 115.800 51.600 120.400 ;
        RECT 58.800 116.200 59.600 120.400 ;
        RECT 62.000 115.800 62.800 120.400 ;
        RECT 63.600 115.800 64.400 120.400 ;
        RECT 66.800 112.200 67.600 120.400 ;
        RECT 70.000 115.800 70.800 120.400 ;
        RECT 73.200 115.800 74.000 120.400 ;
        RECT 74.800 111.800 75.600 120.400 ;
        RECT 79.600 115.800 80.400 120.400 ;
        RECT 82.800 115.800 83.600 120.400 ;
        RECT 85.000 115.800 85.800 120.400 ;
        RECT 89.200 111.800 90.000 120.400 ;
        RECT 94.000 113.000 94.800 120.400 ;
        RECT 98.800 115.800 99.600 120.400 ;
        RECT 102.000 111.800 102.800 120.400 ;
        RECT 107.600 115.800 108.400 120.400 ;
        RECT 110.800 115.800 111.600 120.400 ;
        RECT 116.400 112.000 117.200 120.400 ;
        RECT 122.800 111.800 123.600 120.400 ;
        RECT 126.000 112.000 126.800 120.400 ;
        RECT 131.600 115.800 132.400 120.400 ;
        RECT 134.800 115.800 135.600 120.400 ;
        RECT 140.400 111.800 141.200 120.400 ;
        RECT 149.000 115.800 149.800 120.400 ;
        RECT 153.200 111.800 154.000 120.400 ;
        RECT 154.800 111.800 155.600 120.400 ;
        RECT 159.000 115.800 159.800 120.400 ;
        RECT 162.800 115.800 163.600 120.400 ;
        RECT 167.600 111.800 168.400 120.400 ;
        RECT 169.200 115.800 170.000 120.400 ;
        RECT 172.400 116.200 173.200 120.400 ;
        RECT 177.200 113.800 178.000 120.400 ;
        RECT 190.000 113.000 190.800 120.400 ;
        RECT 2.800 81.600 3.600 89.000 ;
        RECT 7.600 81.600 8.400 90.200 ;
        RECT 13.200 81.600 14.000 86.200 ;
        RECT 16.400 81.600 17.200 86.200 ;
        RECT 22.000 81.600 22.800 90.000 ;
        RECT 25.200 81.600 26.000 90.200 ;
        RECT 29.400 81.600 30.200 86.200 ;
        RECT 34.800 81.600 35.600 90.200 ;
        RECT 39.600 81.600 40.400 90.200 ;
        RECT 41.200 81.600 42.000 86.200 ;
        RECT 44.400 81.600 45.200 86.200 ;
        RECT 47.600 81.600 48.400 86.200 ;
        RECT 50.800 81.600 51.600 89.000 ;
        RECT 58.800 81.600 59.600 86.200 ;
        RECT 62.000 81.600 62.800 89.800 ;
        RECT 65.200 81.600 66.000 86.200 ;
        RECT 68.400 81.600 69.200 86.200 ;
        RECT 73.200 81.600 74.000 90.200 ;
        RECT 76.400 81.600 77.200 89.000 ;
        RECT 82.800 81.600 83.600 90.200 ;
        RECT 87.600 81.600 88.400 90.200 ;
        RECT 90.800 81.600 91.600 90.200 ;
        RECT 96.400 81.600 97.200 86.200 ;
        RECT 99.600 81.600 100.400 86.200 ;
        RECT 105.200 81.600 106.000 90.000 ;
        RECT 110.000 81.600 110.800 89.000 ;
        RECT 114.800 81.600 115.600 86.200 ;
        RECT 118.000 81.600 118.800 86.200 ;
        RECT 121.200 81.600 122.000 89.000 ;
        RECT 127.600 81.600 128.400 85.800 ;
        RECT 130.800 81.600 131.600 86.200 ;
        RECT 134.000 81.600 134.800 89.000 ;
        RECT 143.600 81.600 144.400 86.200 ;
        RECT 147.400 81.600 148.200 86.200 ;
        RECT 151.600 81.600 152.400 90.200 ;
        RECT 156.400 81.600 157.200 89.000 ;
        RECT 159.600 81.600 160.400 86.200 ;
        RECT 164.400 81.600 165.200 88.200 ;
        RECT 177.200 81.600 178.000 89.000 ;
        RECT 182.000 81.600 182.800 86.200 ;
        RECT 185.200 81.600 186.000 89.000 ;
        RECT 190.000 81.600 190.800 89.000 ;
        RECT 0.400 80.400 194.800 81.600 ;
        RECT 2.800 73.000 3.600 80.400 ;
        RECT 7.600 76.200 8.400 80.400 ;
        RECT 10.800 75.800 11.600 80.400 ;
        RECT 12.400 71.800 13.200 80.400 ;
        RECT 16.600 75.800 17.400 80.400 ;
        RECT 22.000 71.800 22.800 80.400 ;
        RECT 23.600 75.800 24.400 80.400 ;
        RECT 26.800 75.800 27.600 80.400 ;
        RECT 28.400 75.800 29.200 80.400 ;
        RECT 31.600 71.800 32.400 80.400 ;
        RECT 35.800 75.800 36.600 80.400 ;
        RECT 41.200 71.800 42.000 80.400 ;
        RECT 44.400 72.000 45.200 80.400 ;
        RECT 50.000 75.800 50.800 80.400 ;
        RECT 53.200 75.800 54.000 80.400 ;
        RECT 58.800 71.800 59.600 80.400 ;
        RECT 66.800 75.800 67.600 80.400 ;
        RECT 71.600 73.000 72.400 80.400 ;
        RECT 74.800 71.800 75.600 80.400 ;
        RECT 78.000 71.800 78.800 80.400 ;
        RECT 81.200 71.800 82.000 80.400 ;
        RECT 84.400 71.800 85.200 80.400 ;
        RECT 87.600 71.800 88.400 80.400 ;
        RECT 90.800 73.000 91.600 80.400 ;
        RECT 94.600 75.800 95.400 80.400 ;
        RECT 98.800 71.800 99.600 80.400 ;
        RECT 103.600 73.000 104.400 80.400 ;
        RECT 108.400 72.000 109.200 80.400 ;
        RECT 114.000 75.800 114.800 80.400 ;
        RECT 117.200 75.800 118.000 80.400 ;
        RECT 122.800 71.800 123.600 80.400 ;
        RECT 126.000 75.800 126.800 80.400 ;
        RECT 129.200 71.800 130.000 80.400 ;
        RECT 133.400 75.800 134.200 80.400 ;
        RECT 140.400 75.800 141.200 80.400 ;
        RECT 143.600 72.200 144.400 80.400 ;
        RECT 148.400 75.800 149.200 80.400 ;
        RECT 150.000 75.800 150.800 80.400 ;
        RECT 153.200 75.800 154.000 80.400 ;
        RECT 156.400 71.800 157.200 80.400 ;
        RECT 162.000 75.800 162.800 80.400 ;
        RECT 165.200 75.800 166.000 80.400 ;
        RECT 170.800 72.000 171.600 80.400 ;
        RECT 175.600 72.000 176.400 80.400 ;
        RECT 181.200 75.800 182.000 80.400 ;
        RECT 184.400 75.800 185.200 80.400 ;
        RECT 190.000 71.800 190.800 80.400 ;
        RECT 2.800 41.600 3.600 49.000 ;
        RECT 7.600 41.600 8.400 50.200 ;
        RECT 13.200 41.600 14.000 46.200 ;
        RECT 16.400 41.600 17.200 46.200 ;
        RECT 22.000 41.600 22.800 50.000 ;
        RECT 25.200 41.600 26.000 46.200 ;
        RECT 28.400 41.600 29.200 49.800 ;
        RECT 31.600 41.600 32.400 50.200 ;
        RECT 34.800 41.600 35.600 50.200 ;
        RECT 38.000 41.600 38.800 50.200 ;
        RECT 41.200 41.600 42.000 50.200 ;
        RECT 44.400 41.600 45.200 50.200 ;
        RECT 52.400 41.600 53.200 50.000 ;
        RECT 58.000 41.600 58.800 46.200 ;
        RECT 61.200 41.600 62.000 46.200 ;
        RECT 66.800 41.600 67.600 50.200 ;
        RECT 70.000 41.600 70.800 46.200 ;
        RECT 73.200 41.600 74.000 46.200 ;
        RECT 74.800 41.600 75.600 50.200 ;
        RECT 82.800 41.600 83.600 49.000 ;
        RECT 86.000 41.600 86.800 46.200 ;
        RECT 89.200 41.600 90.000 46.200 ;
        RECT 90.800 41.600 91.600 50.200 ;
        RECT 94.000 41.600 94.800 50.200 ;
        RECT 97.200 41.600 98.000 50.200 ;
        RECT 100.400 41.600 101.200 50.200 ;
        RECT 103.600 41.600 104.400 50.200 ;
        RECT 105.200 41.600 106.000 46.200 ;
        RECT 108.400 41.600 109.200 46.200 ;
        RECT 110.000 41.600 110.800 50.200 ;
        RECT 124.400 41.600 125.200 48.200 ;
        RECT 127.600 41.600 128.400 50.200 ;
        RECT 131.800 41.600 132.600 46.200 ;
        RECT 140.400 41.600 141.200 49.800 ;
        RECT 143.600 41.600 144.400 46.200 ;
        RECT 145.200 41.600 146.000 46.200 ;
        RECT 148.400 41.600 149.200 46.200 ;
        RECT 150.000 41.600 150.800 46.200 ;
        RECT 153.200 41.600 154.000 49.800 ;
        RECT 156.400 41.600 157.200 46.200 ;
        RECT 159.600 41.600 160.400 45.800 ;
        RECT 164.400 41.600 165.200 45.800 ;
        RECT 167.600 41.600 168.400 46.200 ;
        RECT 169.200 41.600 170.000 50.200 ;
        RECT 175.600 41.600 176.400 49.800 ;
        RECT 178.800 41.600 179.600 46.200 ;
        RECT 180.400 41.600 181.200 46.200 ;
        RECT 183.600 41.600 184.400 46.200 ;
        RECT 186.800 41.600 187.600 49.000 ;
        RECT 191.600 41.600 192.400 49.000 ;
        RECT 0.400 40.400 194.800 41.600 ;
        RECT 2.800 31.800 3.600 40.400 ;
        RECT 8.400 35.800 9.200 40.400 ;
        RECT 11.600 35.800 12.400 40.400 ;
        RECT 17.200 32.000 18.000 40.400 ;
        RECT 21.000 35.800 21.800 40.400 ;
        RECT 25.200 31.800 26.000 40.400 ;
        RECT 26.800 31.800 27.600 40.400 ;
        RECT 32.200 35.800 33.000 40.400 ;
        RECT 36.400 31.800 37.200 40.400 ;
        RECT 38.000 35.800 38.800 40.400 ;
        RECT 41.200 35.800 42.000 40.400 ;
        RECT 43.400 35.800 44.200 40.400 ;
        RECT 47.600 31.800 48.400 40.400 ;
        RECT 49.200 31.800 50.000 40.400 ;
        RECT 58.800 35.800 59.600 40.400 ;
        RECT 62.000 35.800 62.800 40.400 ;
        RECT 63.600 35.800 64.400 40.400 ;
        RECT 66.800 32.200 67.600 40.400 ;
        RECT 71.600 36.200 72.400 40.400 ;
        RECT 74.800 35.800 75.600 40.400 ;
        RECT 78.000 32.200 78.800 40.400 ;
        RECT 81.200 35.800 82.000 40.400 ;
        RECT 84.400 33.000 85.200 40.400 ;
        RECT 89.200 31.800 90.000 40.400 ;
        RECT 93.400 35.800 94.200 40.400 ;
        RECT 96.200 35.800 97.000 40.400 ;
        RECT 100.400 31.800 101.200 40.400 ;
        RECT 103.600 33.000 104.400 40.400 ;
        RECT 110.000 35.800 110.800 40.400 ;
        RECT 111.600 31.800 112.400 40.400 ;
        RECT 115.800 35.800 116.600 40.400 ;
        RECT 118.000 31.800 118.800 40.400 ;
        RECT 122.200 35.800 123.000 40.400 ;
        RECT 127.600 31.800 128.400 40.400 ;
        RECT 135.600 32.000 136.400 40.400 ;
        RECT 141.200 35.800 142.000 40.400 ;
        RECT 144.400 35.800 145.200 40.400 ;
        RECT 150.000 31.800 150.800 40.400 ;
        RECT 154.800 31.800 155.600 40.400 ;
        RECT 160.400 35.800 161.200 40.400 ;
        RECT 163.600 35.800 164.400 40.400 ;
        RECT 169.200 32.000 170.000 40.400 ;
        RECT 174.000 32.000 174.800 40.400 ;
        RECT 179.600 35.800 180.400 40.400 ;
        RECT 182.800 35.800 183.600 40.400 ;
        RECT 188.400 31.800 189.200 40.400 ;
        RECT 2.800 1.600 3.600 9.000 ;
        RECT 7.600 1.600 8.400 10.200 ;
        RECT 13.200 1.600 14.000 6.200 ;
        RECT 16.400 1.600 17.200 6.200 ;
        RECT 22.000 1.600 22.800 10.000 ;
        RECT 28.400 1.600 29.200 9.000 ;
        RECT 33.200 1.600 34.000 9.800 ;
        RECT 36.400 1.600 37.200 6.200 ;
        RECT 39.600 1.600 40.400 9.000 ;
        RECT 47.600 1.600 48.400 10.200 ;
        RECT 55.600 1.600 56.400 10.000 ;
        RECT 61.200 1.600 62.000 6.200 ;
        RECT 64.400 1.600 65.200 6.200 ;
        RECT 70.000 1.600 70.800 10.200 ;
        RECT 74.800 1.600 75.600 9.000 ;
        RECT 79.600 1.600 80.400 9.000 ;
        RECT 84.400 1.600 85.200 9.000 ;
        RECT 89.200 1.600 90.000 9.000 ;
        RECT 94.000 1.600 94.800 9.000 ;
        RECT 98.800 1.600 99.600 10.200 ;
        RECT 104.400 1.600 105.200 6.200 ;
        RECT 107.600 1.600 108.400 6.200 ;
        RECT 113.200 1.600 114.000 10.000 ;
        RECT 116.400 1.600 117.200 6.200 ;
        RECT 119.600 1.600 120.400 6.200 ;
        RECT 122.800 1.600 123.600 10.000 ;
        RECT 128.400 1.600 129.200 6.200 ;
        RECT 131.600 1.600 132.400 6.200 ;
        RECT 137.200 1.600 138.000 10.200 ;
        RECT 146.800 1.600 147.600 9.000 ;
        RECT 151.600 1.600 152.400 9.000 ;
        RECT 156.400 1.600 157.200 9.000 ;
        RECT 161.200 1.600 162.000 9.000 ;
        RECT 164.400 1.600 165.200 6.200 ;
        RECT 169.200 1.600 170.000 9.000 ;
        RECT 176.600 1.600 177.400 10.200 ;
        RECT 182.000 1.600 182.800 9.800 ;
        RECT 185.200 1.600 186.000 6.200 ;
        RECT 190.000 1.600 190.800 9.000 ;
        RECT 0.400 0.400 194.800 1.600 ;
      LAYER via1 ;
        RECT 52.600 160.600 53.400 161.400 ;
        RECT 54.000 160.600 54.800 161.400 ;
        RECT 55.400 160.600 56.200 161.400 ;
        RECT 52.600 120.600 53.400 121.400 ;
        RECT 54.000 120.600 54.800 121.400 ;
        RECT 55.400 120.600 56.200 121.400 ;
        RECT 52.600 80.600 53.400 81.400 ;
        RECT 54.000 80.600 54.800 81.400 ;
        RECT 55.400 80.600 56.200 81.400 ;
        RECT 52.600 40.600 53.400 41.400 ;
        RECT 54.000 40.600 54.800 41.400 ;
        RECT 55.400 40.600 56.200 41.400 ;
        RECT 52.600 0.600 53.400 1.400 ;
        RECT 54.000 0.600 54.800 1.400 ;
        RECT 55.400 0.600 56.200 1.400 ;
      LAYER metal2 ;
        RECT 52.000 160.600 56.800 161.400 ;
        RECT 52.000 120.600 56.800 121.400 ;
        RECT 52.000 80.600 56.800 81.400 ;
        RECT 52.000 40.600 56.800 41.400 ;
        RECT 52.000 0.600 56.800 1.400 ;
      LAYER via2 ;
        RECT 52.600 160.600 53.400 161.400 ;
        RECT 54.000 160.600 54.800 161.400 ;
        RECT 55.400 160.600 56.200 161.400 ;
        RECT 52.600 120.600 53.400 121.400 ;
        RECT 54.000 120.600 54.800 121.400 ;
        RECT 55.400 120.600 56.200 121.400 ;
        RECT 52.600 80.600 53.400 81.400 ;
        RECT 54.000 80.600 54.800 81.400 ;
        RECT 55.400 80.600 56.200 81.400 ;
        RECT 52.600 40.600 53.400 41.400 ;
        RECT 54.000 40.600 54.800 41.400 ;
        RECT 55.400 40.600 56.200 41.400 ;
        RECT 52.600 0.600 53.400 1.400 ;
        RECT 54.000 0.600 54.800 1.400 ;
        RECT 55.400 0.600 56.200 1.400 ;
      LAYER metal3 ;
        RECT 52.000 160.400 56.800 161.600 ;
        RECT 52.000 120.400 56.800 121.600 ;
        RECT 52.000 80.400 56.800 81.600 ;
        RECT 52.000 40.400 56.800 41.600 ;
        RECT 52.000 0.400 56.800 1.600 ;
      LAYER via3 ;
        RECT 52.400 160.600 53.200 161.400 ;
        RECT 54.000 160.600 54.800 161.400 ;
        RECT 55.600 160.600 56.400 161.400 ;
        RECT 52.400 120.600 53.200 121.400 ;
        RECT 54.000 120.600 54.800 121.400 ;
        RECT 55.600 120.600 56.400 121.400 ;
        RECT 52.400 80.600 53.200 81.400 ;
        RECT 54.000 80.600 54.800 81.400 ;
        RECT 55.600 80.600 56.400 81.400 ;
        RECT 52.400 40.600 53.200 41.400 ;
        RECT 54.000 40.600 54.800 41.400 ;
        RECT 55.600 40.600 56.400 41.400 ;
        RECT 52.400 0.600 53.200 1.400 ;
        RECT 54.000 0.600 54.800 1.400 ;
        RECT 55.600 0.600 56.400 1.400 ;
      LAYER metal4 ;
        RECT 52.000 -4.000 56.800 184.000 ;
    END
  END vdd
  PIN gnd
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.400 180.400 194.800 181.600 ;
        RECT 1.200 175.800 2.000 180.400 ;
        RECT 4.400 175.800 5.200 180.400 ;
        RECT 7.600 175.800 8.400 180.400 ;
        RECT 10.800 175.800 11.600 180.400 ;
        RECT 14.000 175.800 14.800 180.400 ;
        RECT 17.200 176.000 18.000 180.400 ;
        RECT 22.800 177.800 23.600 180.400 ;
        RECT 26.000 177.800 27.000 180.400 ;
        RECT 31.600 175.800 32.400 180.400 ;
        RECT 36.400 175.800 37.200 180.400 ;
        RECT 41.200 175.800 42.000 180.400 ;
        RECT 46.600 177.800 47.600 180.400 ;
        RECT 50.000 177.800 50.800 180.400 ;
        RECT 55.600 176.000 56.400 180.400 ;
        RECT 65.200 175.800 66.000 180.400 ;
        RECT 70.000 175.800 70.800 180.400 ;
        RECT 74.800 175.800 75.600 180.400 ;
        RECT 79.600 176.000 80.400 180.400 ;
        RECT 85.200 177.800 86.000 180.400 ;
        RECT 88.400 177.800 89.400 180.400 ;
        RECT 94.000 175.800 94.800 180.400 ;
        RECT 98.800 175.800 99.600 180.400 ;
        RECT 103.600 175.800 104.400 180.400 ;
        RECT 108.400 176.000 109.200 180.400 ;
        RECT 114.000 177.800 114.800 180.400 ;
        RECT 117.200 177.800 118.200 180.400 ;
        RECT 122.800 175.800 123.600 180.400 ;
        RECT 127.600 175.800 128.400 180.400 ;
        RECT 132.400 175.800 133.200 180.400 ;
        RECT 142.000 176.000 142.800 180.400 ;
        RECT 147.600 177.800 148.400 180.400 ;
        RECT 150.800 177.800 151.800 180.400 ;
        RECT 156.400 175.800 157.200 180.400 ;
        RECT 161.200 175.800 162.000 180.400 ;
        RECT 166.000 175.800 166.800 180.400 ;
        RECT 171.400 177.800 172.400 180.400 ;
        RECT 174.800 177.800 175.600 180.400 ;
        RECT 180.400 176.000 181.200 180.400 ;
        RECT 185.200 176.200 186.000 180.400 ;
        RECT 188.400 177.800 189.200 180.400 ;
        RECT 191.600 175.800 192.400 180.400 ;
        RECT 2.800 141.600 3.600 146.000 ;
        RECT 8.400 141.600 9.200 144.200 ;
        RECT 11.600 141.600 12.600 144.200 ;
        RECT 17.200 141.600 18.000 146.200 ;
        RECT 22.000 141.600 22.800 146.000 ;
        RECT 27.600 141.600 28.400 144.200 ;
        RECT 30.800 141.600 31.800 144.200 ;
        RECT 36.400 141.600 37.200 146.200 ;
        RECT 41.800 141.600 42.600 146.000 ;
        RECT 46.000 141.600 46.800 144.200 ;
        RECT 49.800 141.600 50.600 146.200 ;
        RECT 54.000 141.600 54.800 144.200 ;
        RECT 60.400 141.600 61.200 146.200 ;
        RECT 65.200 141.600 66.000 144.200 ;
        RECT 68.400 141.600 69.200 144.200 ;
        RECT 72.600 141.600 73.400 146.200 ;
        RECT 78.000 141.600 78.800 146.200 ;
        RECT 79.600 141.600 80.400 144.200 ;
        RECT 84.400 141.600 85.200 145.800 ;
        RECT 87.600 141.600 88.400 144.200 ;
        RECT 89.800 141.600 90.600 146.200 ;
        RECT 94.000 141.600 94.800 144.200 ;
        RECT 98.200 141.600 99.000 146.000 ;
        RECT 102.000 141.600 102.800 146.200 ;
        RECT 105.200 141.600 106.000 146.200 ;
        RECT 108.400 141.600 109.200 146.200 ;
        RECT 111.600 141.600 112.400 146.200 ;
        RECT 114.800 141.600 115.600 146.200 ;
        RECT 117.000 141.600 117.800 146.200 ;
        RECT 121.200 141.600 122.000 144.200 ;
        RECT 126.000 141.600 126.800 145.400 ;
        RECT 129.200 141.600 130.000 146.200 ;
        RECT 139.400 141.600 140.200 146.200 ;
        RECT 143.600 141.600 144.400 144.200 ;
        RECT 146.800 141.600 147.600 145.400 ;
        RECT 151.600 141.600 152.400 144.200 ;
        RECT 154.800 141.600 155.600 144.200 ;
        RECT 158.000 141.600 158.800 146.000 ;
        RECT 163.600 141.600 164.400 144.200 ;
        RECT 166.800 141.600 167.800 144.200 ;
        RECT 172.400 141.600 173.200 146.200 ;
        RECT 177.200 141.600 178.000 146.200 ;
        RECT 182.600 141.600 183.600 144.200 ;
        RECT 186.000 141.600 186.800 144.200 ;
        RECT 191.600 141.600 192.400 146.000 ;
        RECT 0.400 140.400 194.800 141.600 ;
        RECT 2.800 135.800 3.600 140.400 ;
        RECT 7.600 135.800 8.400 140.400 ;
        RECT 11.400 135.800 12.200 140.400 ;
        RECT 15.600 137.800 16.400 140.400 ;
        RECT 18.800 136.600 19.600 140.400 ;
        RECT 23.600 137.800 24.400 140.400 ;
        RECT 26.800 135.800 27.600 140.400 ;
        RECT 33.200 136.200 34.000 140.400 ;
        RECT 36.400 137.800 37.200 140.400 ;
        RECT 38.600 135.800 39.400 140.400 ;
        RECT 42.800 137.800 43.600 140.400 ;
        RECT 44.400 137.800 45.200 140.400 ;
        RECT 47.600 137.800 48.400 140.400 ;
        RECT 50.800 137.800 51.600 140.400 ;
        RECT 57.800 135.800 58.600 140.400 ;
        RECT 62.000 137.800 62.800 140.400 ;
        RECT 66.800 135.800 67.600 140.400 ;
        RECT 71.600 136.600 72.400 140.400 ;
        RECT 74.800 137.800 75.600 140.400 ;
        RECT 78.000 137.800 78.800 140.400 ;
        RECT 82.800 135.800 83.600 140.400 ;
        RECT 86.000 136.000 86.800 140.400 ;
        RECT 91.600 137.800 92.400 140.400 ;
        RECT 94.800 137.800 95.800 140.400 ;
        RECT 100.400 135.800 101.200 140.400 ;
        RECT 105.200 136.000 106.000 140.400 ;
        RECT 110.800 137.800 111.600 140.400 ;
        RECT 114.000 137.800 115.000 140.400 ;
        RECT 119.600 135.800 120.400 140.400 ;
        RECT 122.800 137.800 123.600 140.400 ;
        RECT 126.000 137.800 126.800 140.400 ;
        RECT 130.800 135.800 131.600 140.400 ;
        RECT 132.400 137.800 133.200 140.400 ;
        RECT 136.600 135.800 137.400 140.400 ;
        RECT 143.600 137.800 144.400 140.400 ;
        RECT 146.800 137.800 147.600 140.400 ;
        RECT 150.000 137.800 150.800 140.400 ;
        RECT 152.200 135.800 153.000 140.400 ;
        RECT 156.400 137.800 157.200 140.400 ;
        RECT 159.600 136.600 160.400 140.400 ;
        RECT 164.400 135.800 165.200 140.400 ;
        RECT 169.200 137.800 170.000 140.400 ;
        RECT 173.400 135.800 174.200 140.400 ;
        RECT 177.200 135.800 178.000 140.400 ;
        RECT 182.600 137.800 183.600 140.400 ;
        RECT 186.000 137.800 186.800 140.400 ;
        RECT 191.600 136.000 192.400 140.400 ;
        RECT 2.800 101.600 3.600 106.200 ;
        RECT 7.600 101.600 8.400 106.000 ;
        RECT 13.200 101.600 14.000 104.200 ;
        RECT 16.400 101.600 17.400 104.200 ;
        RECT 22.000 101.600 22.800 106.200 ;
        RECT 27.400 101.600 28.200 106.000 ;
        RECT 31.600 101.600 32.400 104.200 ;
        RECT 34.800 101.600 35.600 104.200 ;
        RECT 38.000 101.600 38.800 104.200 ;
        RECT 41.200 101.600 42.000 105.400 ;
        RECT 50.800 101.600 51.600 108.200 ;
        RECT 62.000 101.600 62.800 108.200 ;
        RECT 66.200 101.600 67.000 106.000 ;
        RECT 70.000 101.600 70.800 106.200 ;
        RECT 74.800 101.600 75.600 104.200 ;
        RECT 78.000 101.600 78.800 104.200 ;
        RECT 79.600 101.600 80.400 106.200 ;
        RECT 87.600 101.600 88.400 105.400 ;
        RECT 90.800 101.600 91.600 104.200 ;
        RECT 95.000 101.600 95.800 106.200 ;
        RECT 98.800 101.600 99.600 104.200 ;
        RECT 102.000 101.600 102.800 106.000 ;
        RECT 107.600 101.600 108.400 104.200 ;
        RECT 110.800 101.600 111.800 104.200 ;
        RECT 116.400 101.600 117.200 106.200 ;
        RECT 119.600 101.600 120.400 104.200 ;
        RECT 122.800 101.600 123.600 104.200 ;
        RECT 126.000 101.600 126.800 106.200 ;
        RECT 131.400 101.600 132.400 104.200 ;
        RECT 134.800 101.600 135.600 104.200 ;
        RECT 140.400 101.600 141.200 106.000 ;
        RECT 151.600 101.600 152.400 105.400 ;
        RECT 156.400 101.600 157.200 105.400 ;
        RECT 162.800 101.600 163.600 104.200 ;
        RECT 164.400 101.600 165.200 104.200 ;
        RECT 167.600 101.600 168.400 104.200 ;
        RECT 169.200 101.600 170.000 108.200 ;
        RECT 177.200 101.600 178.000 104.200 ;
        RECT 180.400 101.600 181.200 103.800 ;
        RECT 190.000 101.600 190.800 106.200 ;
        RECT 0.400 100.400 194.800 101.600 ;
        RECT 2.800 95.800 3.600 100.400 ;
        RECT 7.600 96.000 8.400 100.400 ;
        RECT 13.200 97.800 14.000 100.400 ;
        RECT 16.400 97.800 17.400 100.400 ;
        RECT 22.000 95.800 22.800 100.400 ;
        RECT 26.800 96.600 27.600 100.400 ;
        RECT 31.600 97.800 32.400 100.400 ;
        RECT 34.800 97.800 35.600 100.400 ;
        RECT 36.400 97.800 37.200 100.400 ;
        RECT 39.600 97.800 40.400 100.400 ;
        RECT 41.200 97.800 42.000 100.400 ;
        RECT 44.400 95.800 45.200 100.400 ;
        RECT 50.800 95.800 51.600 100.400 ;
        RECT 61.400 96.000 62.200 100.400 ;
        RECT 65.200 95.800 66.000 100.400 ;
        RECT 70.000 97.800 70.800 100.400 ;
        RECT 73.200 97.800 74.000 100.400 ;
        RECT 76.400 95.800 77.200 100.400 ;
        RECT 79.600 97.800 80.400 100.400 ;
        RECT 82.800 97.800 83.600 100.400 ;
        RECT 84.400 97.800 85.200 100.400 ;
        RECT 87.600 97.800 88.400 100.400 ;
        RECT 90.800 96.000 91.600 100.400 ;
        RECT 96.400 97.800 97.200 100.400 ;
        RECT 99.600 97.800 100.600 100.400 ;
        RECT 105.200 95.800 106.000 100.400 ;
        RECT 110.000 95.800 110.800 100.400 ;
        RECT 114.800 97.800 115.600 100.400 ;
        RECT 118.000 97.800 118.800 100.400 ;
        RECT 120.200 95.800 121.000 100.400 ;
        RECT 124.400 97.800 125.200 100.400 ;
        RECT 130.800 93.800 131.600 100.400 ;
        RECT 133.000 95.800 133.800 100.400 ;
        RECT 137.200 97.800 138.000 100.400 ;
        RECT 143.600 97.800 144.400 100.400 ;
        RECT 150.000 96.600 150.800 100.400 ;
        RECT 153.200 97.800 154.000 100.400 ;
        RECT 157.400 95.800 158.200 100.400 ;
        RECT 159.600 97.800 160.400 100.400 ;
        RECT 164.400 97.800 165.200 100.400 ;
        RECT 167.600 98.200 168.400 100.400 ;
        RECT 177.200 95.800 178.000 100.400 ;
        RECT 182.000 97.800 182.800 100.400 ;
        RECT 185.200 95.800 186.000 100.400 ;
        RECT 190.000 95.800 190.800 100.400 ;
        RECT 2.800 61.600 3.600 66.200 ;
        RECT 10.800 61.600 11.600 68.200 ;
        RECT 14.000 61.600 14.800 65.400 ;
        RECT 18.800 61.600 19.600 64.200 ;
        RECT 22.000 61.600 22.800 64.200 ;
        RECT 23.600 61.600 24.400 66.200 ;
        RECT 28.400 61.600 29.200 64.200 ;
        RECT 33.200 61.600 34.000 65.400 ;
        RECT 38.000 61.600 38.800 64.200 ;
        RECT 41.200 61.600 42.000 64.200 ;
        RECT 44.400 61.600 45.200 66.200 ;
        RECT 49.800 61.600 50.800 64.200 ;
        RECT 53.200 61.600 54.000 64.200 ;
        RECT 58.800 61.600 59.600 66.000 ;
        RECT 66.800 61.600 67.600 64.200 ;
        RECT 71.600 61.600 72.400 66.200 ;
        RECT 74.800 61.600 75.600 66.200 ;
        RECT 78.000 61.600 78.800 66.200 ;
        RECT 81.200 61.600 82.000 66.200 ;
        RECT 84.400 61.600 85.200 66.200 ;
        RECT 87.600 61.600 88.400 66.200 ;
        RECT 90.800 61.600 91.600 66.200 ;
        RECT 97.200 61.600 98.000 65.400 ;
        RECT 100.400 61.600 101.200 64.200 ;
        RECT 104.600 61.600 105.400 66.200 ;
        RECT 108.400 61.600 109.200 66.200 ;
        RECT 113.800 61.600 114.800 64.200 ;
        RECT 117.200 61.600 118.000 64.200 ;
        RECT 122.800 61.600 123.600 66.000 ;
        RECT 126.000 61.600 126.800 64.200 ;
        RECT 130.800 61.600 131.600 65.400 ;
        RECT 143.000 61.600 143.800 66.000 ;
        RECT 148.400 61.600 149.200 64.200 ;
        RECT 150.000 61.600 150.800 66.200 ;
        RECT 156.400 61.600 157.200 66.000 ;
        RECT 162.000 61.600 162.800 64.200 ;
        RECT 165.200 61.600 166.200 64.200 ;
        RECT 170.800 61.600 171.600 66.200 ;
        RECT 175.600 61.600 176.400 66.200 ;
        RECT 181.000 61.600 182.000 64.200 ;
        RECT 184.400 61.600 185.200 64.200 ;
        RECT 190.000 61.600 190.800 66.000 ;
        RECT 0.400 60.400 194.800 61.600 ;
        RECT 2.800 55.800 3.600 60.400 ;
        RECT 7.600 56.000 8.400 60.400 ;
        RECT 13.200 57.800 14.000 60.400 ;
        RECT 16.400 57.800 17.400 60.400 ;
        RECT 22.000 55.800 22.800 60.400 ;
        RECT 27.800 56.000 28.600 60.400 ;
        RECT 31.600 55.800 32.400 60.400 ;
        RECT 34.800 55.800 35.600 60.400 ;
        RECT 38.000 55.800 38.800 60.400 ;
        RECT 41.200 55.800 42.000 60.400 ;
        RECT 44.400 55.800 45.200 60.400 ;
        RECT 52.400 55.800 53.200 60.400 ;
        RECT 57.800 57.800 58.800 60.400 ;
        RECT 61.200 57.800 62.000 60.400 ;
        RECT 66.800 56.000 67.600 60.400 ;
        RECT 70.000 55.800 70.800 60.400 ;
        RECT 74.800 57.800 75.600 60.400 ;
        RECT 78.000 57.800 78.800 60.400 ;
        RECT 79.600 57.800 80.400 60.400 ;
        RECT 83.800 55.800 84.600 60.400 ;
        RECT 86.000 55.800 86.800 60.400 ;
        RECT 90.800 55.800 91.600 60.400 ;
        RECT 94.000 55.800 94.800 60.400 ;
        RECT 97.200 55.800 98.000 60.400 ;
        RECT 100.400 55.800 101.200 60.400 ;
        RECT 103.600 55.800 104.400 60.400 ;
        RECT 108.400 55.800 109.200 60.400 ;
        RECT 110.000 57.800 110.800 60.400 ;
        RECT 113.200 57.800 114.000 60.400 ;
        RECT 121.200 58.200 122.000 60.400 ;
        RECT 124.400 57.800 125.200 60.400 ;
        RECT 129.200 56.600 130.000 60.400 ;
        RECT 141.000 56.000 141.800 60.400 ;
        RECT 148.400 55.800 149.200 60.400 ;
        RECT 152.600 56.000 153.400 60.400 ;
        RECT 156.400 53.800 157.200 60.400 ;
        RECT 167.600 53.800 168.400 60.400 ;
        RECT 169.200 57.800 170.000 60.400 ;
        RECT 172.400 57.800 173.200 60.400 ;
        RECT 176.200 56.000 177.000 60.400 ;
        RECT 183.600 55.800 184.400 60.400 ;
        RECT 186.800 55.800 187.600 60.400 ;
        RECT 191.600 55.800 192.400 60.400 ;
        RECT 2.800 21.600 3.600 26.000 ;
        RECT 8.400 21.600 9.200 24.200 ;
        RECT 11.600 21.600 12.600 24.200 ;
        RECT 17.200 21.600 18.000 26.200 ;
        RECT 23.600 21.600 24.400 25.400 ;
        RECT 26.800 21.600 27.600 24.200 ;
        RECT 30.000 21.600 30.800 24.200 ;
        RECT 34.800 21.600 35.600 25.400 ;
        RECT 38.000 21.600 38.800 26.200 ;
        RECT 46.000 21.600 46.800 25.400 ;
        RECT 49.200 21.600 50.000 24.200 ;
        RECT 52.400 21.600 53.200 24.200 ;
        RECT 62.000 21.600 62.800 26.200 ;
        RECT 66.200 21.600 67.000 26.000 ;
        RECT 74.800 21.600 75.600 28.200 ;
        RECT 78.600 21.600 79.400 26.000 ;
        RECT 83.400 21.600 84.200 26.200 ;
        RECT 87.600 21.600 88.400 24.200 ;
        RECT 90.800 21.600 91.600 25.400 ;
        RECT 98.800 21.600 99.600 25.400 ;
        RECT 102.600 21.600 103.400 26.200 ;
        RECT 106.800 21.600 107.600 24.200 ;
        RECT 110.000 21.600 110.800 24.200 ;
        RECT 113.200 21.600 114.000 25.400 ;
        RECT 119.600 21.600 120.400 25.400 ;
        RECT 124.400 21.600 125.200 24.200 ;
        RECT 127.600 21.600 128.400 24.200 ;
        RECT 135.600 21.600 136.400 26.200 ;
        RECT 141.000 21.600 142.000 24.200 ;
        RECT 144.400 21.600 145.200 24.200 ;
        RECT 150.000 21.600 150.800 26.000 ;
        RECT 154.800 21.600 155.600 26.000 ;
        RECT 160.400 21.600 161.200 24.200 ;
        RECT 163.600 21.600 164.600 24.200 ;
        RECT 169.200 21.600 170.000 26.200 ;
        RECT 174.000 21.600 174.800 26.200 ;
        RECT 179.400 21.600 180.400 24.200 ;
        RECT 182.800 21.600 183.600 24.200 ;
        RECT 188.400 21.600 189.200 26.000 ;
        RECT 0.400 20.400 194.800 21.600 ;
        RECT 2.800 15.800 3.600 20.400 ;
        RECT 7.600 16.000 8.400 20.400 ;
        RECT 13.200 17.800 14.000 20.400 ;
        RECT 16.400 17.800 17.400 20.400 ;
        RECT 22.000 15.800 22.800 20.400 ;
        RECT 25.200 17.800 26.000 20.400 ;
        RECT 29.400 15.800 30.200 20.400 ;
        RECT 33.800 16.000 34.600 20.400 ;
        RECT 38.600 15.800 39.400 20.400 ;
        RECT 42.800 17.800 43.600 20.400 ;
        RECT 44.400 17.800 45.200 20.400 ;
        RECT 47.600 17.800 48.400 20.400 ;
        RECT 55.600 15.800 56.400 20.400 ;
        RECT 61.000 17.800 62.000 20.400 ;
        RECT 64.400 17.800 65.200 20.400 ;
        RECT 70.000 16.000 70.800 20.400 ;
        RECT 74.800 15.800 75.600 20.400 ;
        RECT 79.600 15.800 80.400 20.400 ;
        RECT 84.400 15.800 85.200 20.400 ;
        RECT 89.200 15.800 90.000 20.400 ;
        RECT 94.000 15.800 94.800 20.400 ;
        RECT 98.800 16.000 99.600 20.400 ;
        RECT 104.400 17.800 105.200 20.400 ;
        RECT 107.600 17.800 108.600 20.400 ;
        RECT 113.200 15.800 114.000 20.400 ;
        RECT 119.600 15.800 120.400 20.400 ;
        RECT 122.800 15.800 123.600 20.400 ;
        RECT 128.200 17.800 129.200 20.400 ;
        RECT 131.600 17.800 132.400 20.400 ;
        RECT 137.200 16.000 138.000 20.400 ;
        RECT 146.800 15.800 147.600 20.400 ;
        RECT 151.600 15.800 152.400 20.400 ;
        RECT 156.400 15.800 157.200 20.400 ;
        RECT 161.200 15.800 162.000 20.400 ;
        RECT 164.400 17.800 165.200 20.400 ;
        RECT 168.200 15.800 169.000 20.400 ;
        RECT 172.400 17.800 173.200 20.400 ;
        RECT 174.000 17.800 174.800 20.400 ;
        RECT 177.200 16.200 178.000 20.400 ;
        RECT 182.600 16.000 183.400 20.400 ;
        RECT 186.800 17.800 187.600 20.400 ;
        RECT 191.000 15.800 191.800 20.400 ;
      LAYER via1 ;
        RECT 135.800 180.600 136.600 181.400 ;
        RECT 137.200 180.600 138.000 181.400 ;
        RECT 138.600 180.600 139.400 181.400 ;
        RECT 135.800 140.600 136.600 141.400 ;
        RECT 137.200 140.600 138.000 141.400 ;
        RECT 138.600 140.600 139.400 141.400 ;
        RECT 135.800 100.600 136.600 101.400 ;
        RECT 137.200 100.600 138.000 101.400 ;
        RECT 138.600 100.600 139.400 101.400 ;
        RECT 135.800 60.600 136.600 61.400 ;
        RECT 137.200 60.600 138.000 61.400 ;
        RECT 138.600 60.600 139.400 61.400 ;
        RECT 135.800 20.600 136.600 21.400 ;
        RECT 137.200 20.600 138.000 21.400 ;
        RECT 138.600 20.600 139.400 21.400 ;
      LAYER metal2 ;
        RECT 135.200 180.600 140.000 181.400 ;
        RECT 135.200 140.600 140.000 141.400 ;
        RECT 135.200 100.600 140.000 101.400 ;
        RECT 135.200 60.600 140.000 61.400 ;
        RECT 135.200 20.600 140.000 21.400 ;
      LAYER via2 ;
        RECT 135.800 180.600 136.600 181.400 ;
        RECT 137.200 180.600 138.000 181.400 ;
        RECT 138.600 180.600 139.400 181.400 ;
        RECT 135.800 140.600 136.600 141.400 ;
        RECT 137.200 140.600 138.000 141.400 ;
        RECT 138.600 140.600 139.400 141.400 ;
        RECT 135.800 100.600 136.600 101.400 ;
        RECT 137.200 100.600 138.000 101.400 ;
        RECT 138.600 100.600 139.400 101.400 ;
        RECT 135.800 60.600 136.600 61.400 ;
        RECT 137.200 60.600 138.000 61.400 ;
        RECT 138.600 60.600 139.400 61.400 ;
        RECT 135.800 20.600 136.600 21.400 ;
        RECT 137.200 20.600 138.000 21.400 ;
        RECT 138.600 20.600 139.400 21.400 ;
      LAYER metal3 ;
        RECT 135.200 180.400 140.000 181.600 ;
        RECT 135.200 140.400 140.000 141.600 ;
        RECT 135.200 100.400 140.000 101.600 ;
        RECT 135.200 60.400 140.000 61.600 ;
        RECT 135.200 20.400 140.000 21.600 ;
      LAYER via3 ;
        RECT 135.600 180.600 136.400 181.400 ;
        RECT 137.200 180.600 138.000 181.400 ;
        RECT 138.800 180.600 139.600 181.400 ;
        RECT 135.600 140.600 136.400 141.400 ;
        RECT 137.200 140.600 138.000 141.400 ;
        RECT 138.800 140.600 139.600 141.400 ;
        RECT 135.600 100.600 136.400 101.400 ;
        RECT 137.200 100.600 138.000 101.400 ;
        RECT 138.800 100.600 139.600 101.400 ;
        RECT 135.600 60.600 136.400 61.400 ;
        RECT 137.200 60.600 138.000 61.400 ;
        RECT 138.800 60.600 139.600 61.400 ;
        RECT 135.600 20.600 136.400 21.400 ;
        RECT 137.200 20.600 138.000 21.400 ;
        RECT 138.800 20.600 139.600 21.400 ;
      LAYER metal4 ;
        RECT 135.200 -4.000 140.000 184.000 ;
    END
  END gnd
  PIN address_enable
    PORT
      LAYER metal1 ;
        RECT 31.600 104.800 32.400 106.400 ;
        RECT 65.200 93.600 66.000 95.200 ;
        RECT 12.400 68.200 13.200 68.400 ;
        RECT 12.400 67.600 14.000 68.200 ;
        RECT 13.200 67.200 14.000 67.600 ;
        RECT 25.200 52.800 26.000 54.400 ;
        RECT 41.200 31.600 42.000 33.200 ;
        RECT 34.800 28.800 35.600 30.400 ;
        RECT 34.400 13.200 35.600 14.000 ;
        RECT 34.800 12.400 35.400 13.200 ;
        RECT 34.800 11.600 35.600 12.400 ;
      LAYER via1 ;
        RECT 31.600 105.600 32.400 106.400 ;
        RECT 25.200 53.600 26.000 54.400 ;
        RECT 34.800 29.600 35.600 30.400 ;
        RECT 34.800 13.200 35.600 14.000 ;
      LAYER metal2 ;
        RECT 28.400 105.600 29.200 106.400 ;
        RECT 31.600 105.600 32.400 106.400 ;
        RECT 28.500 100.400 29.100 105.600 ;
        RECT 28.400 99.600 29.200 100.400 ;
        RECT 65.200 99.600 66.000 100.400 ;
        RECT 12.400 67.600 13.200 68.400 ;
        RECT 12.500 56.400 13.100 67.600 ;
        RECT 28.500 56.400 29.100 99.600 ;
        RECT 65.300 94.400 65.900 99.600 ;
        RECT 65.200 93.600 66.000 94.400 ;
        RECT 12.400 55.600 13.200 56.400 ;
        RECT 25.200 55.600 26.000 56.400 ;
        RECT 28.400 55.600 29.200 56.400 ;
        RECT 25.300 54.400 25.900 55.600 ;
        RECT 25.200 53.600 26.000 54.400 ;
        RECT 25.300 32.400 25.900 53.600 ;
        RECT 25.200 31.600 26.000 32.400 ;
        RECT 34.800 31.600 35.600 32.400 ;
        RECT 41.200 31.600 42.000 32.400 ;
        RECT 34.900 30.400 35.500 31.600 ;
        RECT 34.800 29.600 35.600 30.400 ;
        RECT 34.900 14.000 35.500 29.600 ;
        RECT 34.800 13.200 35.600 14.000 ;
        RECT 34.900 -1.700 35.500 13.200 ;
        RECT 33.300 -2.300 35.500 -1.700 ;
      LAYER metal3 ;
        RECT 28.400 106.300 29.200 106.400 ;
        RECT 31.600 106.300 32.400 106.400 ;
        RECT 28.400 105.700 32.400 106.300 ;
        RECT 28.400 105.600 29.200 105.700 ;
        RECT 31.600 105.600 32.400 105.700 ;
        RECT 28.400 100.300 29.200 100.400 ;
        RECT 65.200 100.300 66.000 100.400 ;
        RECT 28.400 99.700 66.000 100.300 ;
        RECT 28.400 99.600 29.200 99.700 ;
        RECT 65.200 99.600 66.000 99.700 ;
        RECT 12.400 56.300 13.200 56.400 ;
        RECT 25.200 56.300 26.000 56.400 ;
        RECT 28.400 56.300 29.200 56.400 ;
        RECT 12.400 55.700 29.200 56.300 ;
        RECT 12.400 55.600 13.200 55.700 ;
        RECT 25.200 55.600 26.000 55.700 ;
        RECT 28.400 55.600 29.200 55.700 ;
        RECT 25.200 32.300 26.000 32.400 ;
        RECT 34.800 32.300 35.600 32.400 ;
        RECT 41.200 32.300 42.000 32.400 ;
        RECT 25.200 31.700 42.000 32.300 ;
        RECT 25.200 31.600 26.000 31.700 ;
        RECT 34.800 31.600 35.600 31.700 ;
        RECT 41.200 31.600 42.000 31.700 ;
    END
  END address_enable
  PIN clock
    PORT
      LAYER metal1 ;
        RECT 1.200 173.800 2.000 174.400 ;
        RECT 1.200 173.000 3.000 173.800 ;
        RECT 102.000 148.200 103.800 149.000 ;
        RECT 102.000 147.600 102.800 148.200 ;
        RECT 74.800 68.200 76.600 69.000 ;
        RECT 74.800 67.600 75.600 68.200 ;
        RECT 44.400 53.800 45.200 54.400 ;
        RECT 43.400 53.000 45.200 53.800 ;
        RECT 90.800 53.800 91.600 54.400 ;
        RECT 90.800 53.000 92.600 53.800 ;
      LAYER via1 ;
        RECT 1.200 173.600 2.000 174.400 ;
        RECT 44.400 53.600 45.200 54.400 ;
        RECT 90.800 53.600 91.600 54.400 ;
      LAYER metal2 ;
        RECT 1.200 173.600 2.000 174.400 ;
        RECT 1.300 170.400 1.900 173.600 ;
        RECT 1.200 169.600 2.000 170.400 ;
        RECT 102.000 167.600 102.800 168.400 ;
        RECT 102.100 148.400 102.700 167.600 ;
        RECT 102.000 147.600 102.800 148.400 ;
        RECT 102.100 146.400 102.700 147.600 ;
        RECT 97.200 145.600 98.000 146.400 ;
        RECT 102.000 145.600 102.800 146.400 ;
        RECT 97.300 104.400 97.900 145.600 ;
        RECT 90.800 103.600 91.600 104.400 ;
        RECT 97.200 103.600 98.000 104.400 ;
        RECT 74.800 67.600 75.600 68.400 ;
        RECT 74.900 56.400 75.500 67.600 ;
        RECT 44.400 55.600 45.200 56.400 ;
        RECT 74.800 55.600 75.600 56.400 ;
        RECT 44.500 54.400 45.100 55.600 ;
        RECT 74.900 54.400 75.500 55.600 ;
        RECT 90.900 54.400 91.500 103.600 ;
        RECT 44.400 53.600 45.200 54.400 ;
        RECT 74.800 53.600 75.600 54.400 ;
        RECT 90.800 53.600 91.600 54.400 ;
      LAYER metal3 ;
        RECT 1.200 170.300 2.000 170.400 ;
        RECT -1.900 169.700 2.000 170.300 ;
        RECT 1.200 169.600 2.000 169.700 ;
        RECT 1.300 168.300 1.900 169.600 ;
        RECT 102.000 168.300 102.800 168.400 ;
        RECT 1.300 167.700 102.800 168.300 ;
        RECT 102.000 167.600 102.800 167.700 ;
        RECT 97.200 146.300 98.000 146.400 ;
        RECT 102.000 146.300 102.800 146.400 ;
        RECT 97.200 145.700 102.800 146.300 ;
        RECT 97.200 145.600 98.000 145.700 ;
        RECT 102.000 145.600 102.800 145.700 ;
        RECT 90.800 104.300 91.600 104.400 ;
        RECT 97.200 104.300 98.000 104.400 ;
        RECT 90.800 103.700 98.000 104.300 ;
        RECT 90.800 103.600 91.600 103.700 ;
        RECT 97.200 103.600 98.000 103.700 ;
        RECT 44.400 56.300 45.200 56.400 ;
        RECT 74.800 56.300 75.600 56.400 ;
        RECT 44.400 55.700 75.600 56.300 ;
        RECT 44.400 55.600 45.200 55.700 ;
        RECT 74.800 55.600 75.600 55.700 ;
        RECT 74.800 54.300 75.600 54.400 ;
        RECT 90.800 54.300 91.600 54.400 ;
        RECT 74.800 53.700 91.600 54.300 ;
        RECT 74.800 53.600 75.600 53.700 ;
        RECT 90.800 53.600 91.600 53.700 ;
    END
  END clock
  PIN reset
    PORT
      LAYER metal1 ;
        RECT 188.400 175.600 189.200 177.200 ;
        RECT 94.000 145.600 94.800 146.400 ;
        RECT 93.800 144.800 94.600 145.600 ;
        RECT 42.600 136.400 43.400 137.200 ;
        RECT 42.800 135.600 43.600 136.400 ;
        RECT 177.200 105.600 179.000 106.400 ;
        RECT 62.000 66.300 62.800 66.400 ;
        RECT 66.800 66.300 67.600 66.400 ;
        RECT 62.000 65.700 67.600 66.300 ;
        RECT 62.000 65.600 62.800 65.700 ;
        RECT 66.800 64.800 67.600 65.700 ;
        RECT 127.600 24.800 128.400 26.400 ;
        RECT 172.200 16.400 173.000 17.200 ;
        RECT 172.400 15.600 173.200 16.400 ;
      LAYER via1 ;
        RECT 127.600 25.600 128.400 26.400 ;
      LAYER metal2 ;
        RECT 185.300 176.400 185.900 184.300 ;
        RECT 185.200 175.600 186.000 176.400 ;
        RECT 188.400 175.600 189.200 176.400 ;
        RECT 94.000 145.600 94.800 146.400 ;
        RECT 42.800 135.600 43.600 136.400 ;
        RECT 42.900 116.400 43.500 135.600 ;
        RECT 94.100 116.400 94.700 145.600 ;
        RECT 185.300 126.400 185.900 175.600 ;
        RECT 177.200 125.600 178.000 126.400 ;
        RECT 185.200 125.600 186.000 126.400 ;
        RECT 177.300 116.400 177.900 125.600 ;
        RECT 42.800 115.600 43.600 116.400 ;
        RECT 62.000 115.600 62.800 116.400 ;
        RECT 94.000 115.600 94.800 116.400 ;
        RECT 177.200 115.600 178.000 116.400 ;
        RECT 62.100 66.400 62.700 115.600 ;
        RECT 177.300 106.400 177.900 115.600 ;
        RECT 177.200 105.600 178.000 106.400 ;
        RECT 62.000 65.600 62.800 66.400 ;
        RECT 127.600 25.600 128.400 26.400 ;
        RECT 172.400 23.600 173.200 24.400 ;
        RECT 172.500 16.400 173.100 23.600 ;
        RECT 172.400 15.600 173.200 16.400 ;
      LAYER metal3 ;
        RECT 185.200 176.300 186.000 176.400 ;
        RECT 188.400 176.300 189.200 176.400 ;
        RECT 185.200 175.700 189.200 176.300 ;
        RECT 185.200 175.600 186.000 175.700 ;
        RECT 188.400 175.600 189.200 175.700 ;
        RECT 177.200 126.300 178.000 126.400 ;
        RECT 185.200 126.300 186.000 126.400 ;
        RECT 177.200 125.700 186.000 126.300 ;
        RECT 177.200 125.600 178.000 125.700 ;
        RECT 185.200 125.600 186.000 125.700 ;
        RECT 42.800 116.300 43.600 116.400 ;
        RECT 62.000 116.300 62.800 116.400 ;
        RECT 94.000 116.300 94.800 116.400 ;
        RECT 119.600 116.300 120.400 116.400 ;
        RECT 177.200 116.300 178.000 116.400 ;
        RECT 42.800 115.700 178.000 116.300 ;
        RECT 42.800 115.600 43.600 115.700 ;
        RECT 62.000 115.600 62.800 115.700 ;
        RECT 94.000 115.600 94.800 115.700 ;
        RECT 119.600 115.600 120.400 115.700 ;
        RECT 177.200 115.600 178.000 115.700 ;
        RECT 119.600 26.300 120.400 26.400 ;
        RECT 127.600 26.300 128.400 26.400 ;
        RECT 119.600 25.700 128.400 26.300 ;
        RECT 119.600 25.600 120.400 25.700 ;
        RECT 127.600 25.600 128.400 25.700 ;
        RECT 127.700 24.300 128.300 25.600 ;
        RECT 172.400 24.300 173.200 24.400 ;
        RECT 127.700 23.700 173.200 24.300 ;
        RECT 172.400 23.600 173.200 23.700 ;
      LAYER metal4 ;
        RECT 119.400 25.400 120.600 116.600 ;
    END
  END reset
  PIN address_a[0]
    PORT
      LAYER metal1 ;
        RECT 1.200 111.800 2.000 119.800 ;
        RECT 1.200 109.600 1.800 111.800 ;
        RECT 1.200 102.200 2.000 109.600 ;
      LAYER via1 ;
        RECT 1.200 107.600 2.000 108.400 ;
      LAYER metal2 ;
        RECT 1.200 109.600 2.000 110.400 ;
        RECT 1.300 108.400 1.900 109.600 ;
        RECT 1.200 107.600 2.000 108.400 ;
      LAYER metal3 ;
        RECT 1.200 110.300 2.000 110.400 ;
        RECT -1.900 109.700 2.000 110.300 ;
        RECT 1.200 109.600 2.000 109.700 ;
    END
  END address_a[0]
  PIN address_a[1]
    PORT
      LAYER metal1 ;
        RECT 1.200 52.400 2.000 59.800 ;
        RECT 1.200 50.200 1.800 52.400 ;
        RECT 1.200 42.200 2.000 50.200 ;
      LAYER via1 ;
        RECT 1.200 47.600 2.000 48.400 ;
      LAYER metal2 ;
        RECT 1.200 49.600 2.000 50.400 ;
        RECT 1.300 48.400 1.900 49.600 ;
        RECT 1.200 47.600 2.000 48.400 ;
      LAYER metal3 ;
        RECT 1.200 50.300 2.000 50.400 ;
        RECT -1.900 49.700 2.000 50.300 ;
        RECT 1.200 49.600 2.000 49.700 ;
    END
  END address_a[1]
  PIN address_a[2]
    PORT
      LAYER metal1 ;
        RECT 1.200 71.800 2.000 79.800 ;
        RECT 1.200 69.600 1.800 71.800 ;
        RECT 1.200 62.200 2.000 69.600 ;
      LAYER via1 ;
        RECT 1.200 67.600 2.000 68.400 ;
      LAYER metal2 ;
        RECT 1.200 69.600 2.000 70.400 ;
        RECT 1.300 68.400 1.900 69.600 ;
        RECT 1.200 67.600 2.000 68.400 ;
      LAYER metal3 ;
        RECT 1.200 70.300 2.000 70.400 ;
        RECT -1.900 69.700 2.000 70.300 ;
        RECT 1.200 69.600 2.000 69.700 ;
    END
  END address_a[2]
  PIN address_a[3]
    PORT
      LAYER metal1 ;
        RECT 1.200 92.400 2.000 99.800 ;
        RECT 1.200 90.200 1.800 92.400 ;
        RECT 1.200 82.200 2.000 90.200 ;
      LAYER via1 ;
        RECT 1.200 87.600 2.000 88.400 ;
      LAYER metal2 ;
        RECT 1.200 89.600 2.000 90.400 ;
        RECT 1.300 88.400 1.900 89.600 ;
        RECT 1.200 87.600 2.000 88.400 ;
      LAYER metal3 ;
        RECT 1.200 90.300 2.000 90.400 ;
        RECT -1.900 89.700 2.000 90.300 ;
        RECT 1.200 89.600 2.000 89.700 ;
    END
  END address_a[3]
  PIN address_a[4]
    PORT
      LAYER metal1 ;
        RECT 129.200 172.400 130.000 179.800 ;
        RECT 129.400 170.200 130.000 172.400 ;
        RECT 129.200 162.200 130.000 170.200 ;
      LAYER via1 ;
        RECT 129.200 177.600 130.000 178.400 ;
      LAYER metal2 ;
        RECT 127.700 183.700 129.900 184.300 ;
        RECT 129.300 178.400 129.900 183.700 ;
        RECT 129.200 177.600 130.000 178.400 ;
    END
  END address_a[4]
  PIN address_a[5]
    PORT
      LAYER metal1 ;
        RECT 162.800 172.400 163.600 179.800 ;
        RECT 163.000 170.200 163.600 172.400 ;
        RECT 162.800 162.200 163.600 170.200 ;
      LAYER via1 ;
        RECT 162.800 177.600 163.600 178.400 ;
      LAYER metal2 ;
        RECT 161.300 183.700 163.500 184.300 ;
        RECT 162.900 178.400 163.500 183.700 ;
        RECT 162.800 177.600 163.600 178.400 ;
    END
  END address_a[5]
  PIN address_a[6]
    PORT
      LAYER metal1 ;
        RECT 134.000 172.400 134.800 179.800 ;
        RECT 134.200 170.200 134.800 172.400 ;
        RECT 134.000 162.200 134.800 170.200 ;
      LAYER via1 ;
        RECT 134.000 177.600 134.800 178.400 ;
      LAYER metal2 ;
        RECT 132.500 178.300 133.100 184.300 ;
        RECT 134.000 178.300 134.800 178.400 ;
        RECT 132.500 177.700 134.800 178.300 ;
        RECT 134.000 177.600 134.800 177.700 ;
    END
  END address_a[6]
  PIN address_a[7]
    PORT
      LAYER metal1 ;
        RECT 102.000 172.400 102.800 179.800 ;
        RECT 102.000 170.200 102.600 172.400 ;
        RECT 102.000 162.200 102.800 170.200 ;
      LAYER via1 ;
        RECT 102.000 177.600 102.800 178.400 ;
      LAYER metal2 ;
        RECT 102.100 183.700 104.300 184.300 ;
        RECT 102.100 178.400 102.700 183.700 ;
        RECT 102.000 177.600 102.800 178.400 ;
    END
  END address_a[7]
  PIN address_a[8]
    PORT
      LAYER metal1 ;
        RECT 1.200 132.400 2.000 139.800 ;
        RECT 1.200 130.200 1.800 132.400 ;
        RECT 1.200 122.200 2.000 130.200 ;
      LAYER via1 ;
        RECT 1.200 127.600 2.000 128.400 ;
      LAYER metal2 ;
        RECT 1.200 129.600 2.000 130.400 ;
        RECT 1.300 128.400 1.900 129.600 ;
        RECT 1.200 127.600 2.000 128.400 ;
      LAYER metal3 ;
        RECT 1.200 130.300 2.000 130.400 ;
        RECT -1.900 129.700 2.000 130.300 ;
        RECT 1.200 129.600 2.000 129.700 ;
    END
  END address_a[8]
  PIN address_a[9]
    PORT
      LAYER metal1 ;
        RECT 66.800 172.400 67.600 179.800 ;
        RECT 67.000 170.200 67.600 172.400 ;
        RECT 66.800 162.200 67.600 170.200 ;
      LAYER via1 ;
        RECT 66.800 177.600 67.600 178.400 ;
      LAYER metal2 ;
        RECT 63.700 180.400 64.300 184.300 ;
        RECT 63.600 179.600 64.400 180.400 ;
        RECT 66.800 179.600 67.600 180.400 ;
        RECT 66.900 178.400 67.500 179.600 ;
        RECT 66.800 177.600 67.600 178.400 ;
      LAYER metal3 ;
        RECT 63.600 180.300 64.400 180.400 ;
        RECT 66.800 180.300 67.600 180.400 ;
        RECT 63.600 179.700 67.600 180.300 ;
        RECT 63.600 179.600 64.400 179.700 ;
        RECT 66.800 179.600 67.600 179.700 ;
    END
  END address_a[9]
  PIN address_a[10]
    PORT
      LAYER metal1 ;
        RECT 38.000 172.400 38.800 179.800 ;
        RECT 38.200 170.200 38.800 172.400 ;
        RECT 38.000 162.200 38.800 170.200 ;
      LAYER via1 ;
        RECT 38.000 177.600 38.800 178.400 ;
      LAYER metal2 ;
        RECT 36.500 183.700 38.700 184.300 ;
        RECT 38.100 178.400 38.700 183.700 ;
        RECT 38.000 177.600 38.800 178.400 ;
    END
  END address_a[10]
  PIN address_a[11]
    PORT
      LAYER metal1 ;
        RECT 6.000 132.400 6.800 139.800 ;
        RECT 6.000 130.200 6.600 132.400 ;
        RECT 6.000 122.200 6.800 130.200 ;
      LAYER via1 ;
        RECT 6.000 133.600 6.800 134.400 ;
      LAYER metal2 ;
        RECT 6.000 133.600 6.800 134.400 ;
      LAYER metal3 ;
        RECT 6.000 134.300 6.800 134.400 ;
        RECT -1.900 133.700 6.800 134.300 ;
        RECT 6.000 133.600 6.800 133.700 ;
    END
  END address_a[11]
  PIN address_a[12]
    PORT
      LAYER metal1 ;
        RECT 76.400 172.400 77.200 179.800 ;
        RECT 76.600 170.200 77.200 172.400 ;
        RECT 76.400 162.200 77.200 170.200 ;
      LAYER via1 ;
        RECT 76.400 177.600 77.200 178.400 ;
      LAYER metal2 ;
        RECT 74.900 183.700 77.100 184.300 ;
        RECT 76.500 178.400 77.100 183.700 ;
        RECT 76.400 177.600 77.200 178.400 ;
    END
  END address_a[12]
  PIN address_a[13]
    PORT
      LAYER metal1 ;
        RECT 71.600 172.400 72.400 179.800 ;
        RECT 71.800 170.200 72.400 172.400 ;
        RECT 71.600 162.200 72.400 170.200 ;
      LAYER via1 ;
        RECT 71.600 177.600 72.400 178.400 ;
      LAYER metal2 ;
        RECT 68.500 180.400 69.100 184.300 ;
        RECT 68.400 179.600 69.200 180.400 ;
        RECT 71.600 179.600 72.400 180.400 ;
        RECT 71.700 178.400 72.300 179.600 ;
        RECT 71.600 177.600 72.400 178.400 ;
      LAYER metal3 ;
        RECT 68.400 180.300 69.200 180.400 ;
        RECT 71.600 180.300 72.400 180.400 ;
        RECT 68.400 179.700 72.400 180.300 ;
        RECT 68.400 179.600 69.200 179.700 ;
        RECT 71.600 179.600 72.400 179.700 ;
    END
  END address_a[13]
  PIN address_a[14]
    PORT
      LAYER metal1 ;
        RECT 86.000 12.400 86.800 19.800 ;
        RECT 86.200 10.200 86.800 12.400 ;
        RECT 86.000 2.200 86.800 10.200 ;
      LAYER via1 ;
        RECT 86.000 3.600 86.800 4.400 ;
      LAYER metal2 ;
        RECT 86.000 3.600 86.800 4.400 ;
        RECT 86.100 -1.700 86.700 3.600 ;
        RECT 84.500 -2.300 86.700 -1.700 ;
    END
  END address_a[14]
  PIN address_a[15]
    PORT
      LAYER metal1 ;
        RECT 97.200 172.400 98.000 179.800 ;
        RECT 97.200 170.200 97.800 172.400 ;
        RECT 97.200 162.200 98.000 170.200 ;
      LAYER via1 ;
        RECT 97.200 177.600 98.000 178.400 ;
      LAYER metal2 ;
        RECT 97.300 183.700 99.500 184.300 ;
        RECT 97.300 178.400 97.900 183.700 ;
        RECT 97.200 177.600 98.000 178.400 ;
    END
  END address_a[15]
  PIN address_b[0]
    PORT
      LAYER metal1 ;
        RECT 193.200 172.400 194.000 179.800 ;
        RECT 193.400 170.200 194.000 172.400 ;
        RECT 193.200 162.200 194.000 170.200 ;
      LAYER via1 ;
        RECT 193.200 167.600 194.000 168.400 ;
      LAYER metal2 ;
        RECT 193.200 169.600 194.000 170.400 ;
        RECT 193.300 168.400 193.900 169.600 ;
        RECT 193.200 167.600 194.000 168.400 ;
      LAYER metal3 ;
        RECT 193.200 170.300 194.000 170.400 ;
        RECT 193.200 169.700 197.100 170.300 ;
        RECT 193.200 169.600 194.000 169.700 ;
    END
  END address_b[0]
  PIN address_b[1]
    PORT
      LAYER metal1 ;
        RECT 1.200 12.400 2.000 19.800 ;
        RECT 1.200 10.200 1.800 12.400 ;
        RECT 1.200 2.200 2.000 10.200 ;
      LAYER via1 ;
        RECT 1.200 7.600 2.000 8.400 ;
      LAYER metal2 ;
        RECT 1.200 9.600 2.000 10.400 ;
        RECT 1.300 8.400 1.900 9.600 ;
        RECT 1.200 7.600 2.000 8.400 ;
      LAYER metal3 ;
        RECT 1.200 10.300 2.000 10.400 ;
        RECT -1.900 9.700 2.000 10.300 ;
        RECT 1.200 9.600 2.000 9.700 ;
    END
  END address_b[1]
  PIN address_b[2]
    PORT
      LAYER metal1 ;
        RECT 73.200 12.400 74.000 19.800 ;
        RECT 73.200 10.200 73.800 12.400 ;
        RECT 73.200 2.200 74.000 10.200 ;
      LAYER via1 ;
        RECT 73.200 3.600 74.000 4.400 ;
      LAYER metal2 ;
        RECT 73.200 3.600 74.000 4.400 ;
        RECT 73.300 -2.300 73.900 3.600 ;
    END
  END address_b[2]
  PIN address_b[3]
    PORT
      LAYER metal1 ;
        RECT 81.200 12.400 82.000 19.800 ;
        RECT 81.400 10.200 82.000 12.400 ;
        RECT 81.200 2.200 82.000 10.200 ;
      LAYER via1 ;
        RECT 81.200 3.600 82.000 4.400 ;
      LAYER metal2 ;
        RECT 81.200 3.600 82.000 4.400 ;
        RECT 81.300 -1.700 81.900 3.600 ;
        RECT 79.700 -2.300 81.900 -1.700 ;
    END
  END address_b[3]
  PIN address_b[4]
    PORT
      LAYER metal1 ;
        RECT 95.600 12.400 96.400 19.800 ;
        RECT 95.800 10.200 96.400 12.400 ;
        RECT 95.600 2.200 96.400 10.200 ;
      LAYER via1 ;
        RECT 95.600 3.600 96.400 4.400 ;
      LAYER metal2 ;
        RECT 95.600 3.600 96.400 4.400 ;
        RECT 95.700 -1.700 96.300 3.600 ;
        RECT 94.100 -2.300 96.300 -1.700 ;
    END
  END address_b[4]
  PIN address_b[5]
    PORT
      LAYER metal1 ;
        RECT 90.800 12.400 91.600 19.800 ;
        RECT 91.000 10.200 91.600 12.400 ;
        RECT 90.800 2.200 91.600 10.200 ;
      LAYER via1 ;
        RECT 90.800 3.600 91.600 4.400 ;
      LAYER metal2 ;
        RECT 90.800 3.600 91.600 4.400 ;
        RECT 90.900 -1.700 91.500 3.600 ;
        RECT 89.300 -2.300 91.500 -1.700 ;
    END
  END address_b[5]
  PIN address_b[6]
    PORT
      LAYER metal1 ;
        RECT 148.400 12.400 149.200 19.800 ;
        RECT 148.600 10.200 149.200 12.400 ;
        RECT 148.400 2.200 149.200 10.200 ;
      LAYER via1 ;
        RECT 148.400 3.600 149.200 4.400 ;
      LAYER metal2 ;
        RECT 148.400 3.600 149.200 4.400 ;
        RECT 148.500 2.400 149.100 3.600 ;
        RECT 145.200 1.600 146.000 2.400 ;
        RECT 148.400 1.600 149.200 2.400 ;
        RECT 145.300 -2.300 145.900 1.600 ;
      LAYER metal3 ;
        RECT 145.200 2.300 146.000 2.400 ;
        RECT 148.400 2.300 149.200 2.400 ;
        RECT 145.200 1.700 149.200 2.300 ;
        RECT 145.200 1.600 146.000 1.700 ;
        RECT 148.400 1.600 149.200 1.700 ;
    END
  END address_b[6]
  PIN address_b[7]
    PORT
      LAYER metal1 ;
        RECT 153.200 12.400 154.000 19.800 ;
        RECT 153.400 10.200 154.000 12.400 ;
        RECT 153.200 2.200 154.000 10.200 ;
      LAYER via1 ;
        RECT 153.200 3.600 154.000 4.400 ;
      LAYER metal2 ;
        RECT 153.200 3.600 154.000 4.400 ;
        RECT 153.300 2.400 153.900 3.600 ;
        RECT 150.000 1.600 150.800 2.400 ;
        RECT 153.200 1.600 154.000 2.400 ;
        RECT 150.100 -2.300 150.700 1.600 ;
      LAYER metal3 ;
        RECT 150.000 2.300 150.800 2.400 ;
        RECT 153.200 2.300 154.000 2.400 ;
        RECT 150.000 1.700 154.000 2.300 ;
        RECT 150.000 1.600 150.800 1.700 ;
        RECT 153.200 1.600 154.000 1.700 ;
    END
  END address_b[7]
  PIN address_b[8]
    PORT
      LAYER metal1 ;
        RECT 158.000 12.400 158.800 19.800 ;
        RECT 158.200 10.200 158.800 12.400 ;
        RECT 158.000 2.200 158.800 10.200 ;
      LAYER via1 ;
        RECT 158.000 3.600 158.800 4.400 ;
      LAYER metal2 ;
        RECT 158.000 3.600 158.800 4.400 ;
        RECT 158.100 2.400 158.700 3.600 ;
        RECT 154.800 1.600 155.600 2.400 ;
        RECT 158.000 1.600 158.800 2.400 ;
        RECT 154.900 -2.300 155.500 1.600 ;
      LAYER metal3 ;
        RECT 154.800 2.300 155.600 2.400 ;
        RECT 158.000 2.300 158.800 2.400 ;
        RECT 154.800 1.700 158.800 2.300 ;
        RECT 154.800 1.600 155.600 1.700 ;
        RECT 158.000 1.600 158.800 1.700 ;
    END
  END address_b[8]
  PIN address_b[9]
    PORT
      LAYER metal1 ;
        RECT 162.800 12.400 163.600 19.800 ;
        RECT 163.000 10.200 163.600 12.400 ;
        RECT 162.800 2.200 163.600 10.200 ;
      LAYER via1 ;
        RECT 162.800 3.600 163.600 4.400 ;
      LAYER metal2 ;
        RECT 162.800 3.600 163.600 4.400 ;
        RECT 162.900 -1.700 163.500 3.600 ;
        RECT 161.300 -2.300 163.500 -1.700 ;
    END
  END address_b[9]
  PIN address_b[10]
    PORT
      LAYER metal1 ;
        RECT 193.200 52.400 194.000 59.800 ;
        RECT 193.400 50.200 194.000 52.400 ;
        RECT 193.200 42.200 194.000 50.200 ;
      LAYER via1 ;
        RECT 193.200 47.600 194.000 48.400 ;
      LAYER metal2 ;
        RECT 193.200 49.600 194.000 50.400 ;
        RECT 193.300 48.400 193.900 49.600 ;
        RECT 193.200 47.600 194.000 48.400 ;
      LAYER metal3 ;
        RECT 193.200 50.300 194.000 50.400 ;
        RECT 193.200 49.700 197.100 50.300 ;
        RECT 193.200 49.600 194.000 49.700 ;
    END
  END address_b[10]
  PIN address_b[11]
    PORT
      LAYER metal1 ;
        RECT 188.400 52.400 189.200 59.800 ;
        RECT 188.600 50.200 189.200 52.400 ;
        RECT 188.400 42.200 189.200 50.200 ;
      LAYER via1 ;
        RECT 188.400 53.600 189.200 54.400 ;
      LAYER metal2 ;
        RECT 188.400 53.600 189.200 54.400 ;
      LAYER metal3 ;
        RECT 188.400 54.300 189.200 54.400 ;
        RECT 188.400 53.700 197.100 54.300 ;
        RECT 188.400 53.600 189.200 53.700 ;
    END
  END address_b[11]
  PIN address_b[12]
    PORT
      LAYER metal1 ;
        RECT 186.800 92.400 187.600 99.800 ;
        RECT 187.000 90.200 187.600 92.400 ;
        RECT 186.800 82.200 187.600 90.200 ;
      LAYER via1 ;
        RECT 186.800 87.600 187.600 88.400 ;
      LAYER metal2 ;
        RECT 186.800 89.600 187.600 90.400 ;
        RECT 186.900 88.400 187.500 89.600 ;
        RECT 186.800 87.600 187.600 88.400 ;
      LAYER metal3 ;
        RECT 186.800 90.300 187.600 90.400 ;
        RECT 186.800 89.700 197.100 90.300 ;
        RECT 186.800 89.600 187.600 89.700 ;
    END
  END address_b[12]
  PIN address_b[13]
    PORT
      LAYER metal1 ;
        RECT 191.600 98.300 192.400 99.800 ;
        RECT 193.200 98.300 194.000 98.400 ;
        RECT 191.600 97.700 194.000 98.300 ;
        RECT 191.600 92.400 192.400 97.700 ;
        RECT 193.200 97.600 194.000 97.700 ;
        RECT 191.800 90.200 192.400 92.400 ;
        RECT 191.600 82.200 192.400 90.200 ;
      LAYER metal2 ;
        RECT 193.200 97.600 194.000 98.400 ;
      LAYER metal3 ;
        RECT 193.200 98.300 194.000 98.400 ;
        RECT 193.200 97.700 197.100 98.300 ;
        RECT 193.200 97.600 194.000 97.700 ;
    END
  END address_b[13]
  PIN address_b[14]
    PORT
      LAYER metal1 ;
        RECT 178.800 92.400 179.600 99.800 ;
        RECT 179.000 90.200 179.600 92.400 ;
        RECT 178.800 82.200 179.600 90.200 ;
      LAYER via1 ;
        RECT 178.800 93.600 179.600 94.400 ;
      LAYER metal2 ;
        RECT 178.800 93.600 179.600 94.400 ;
      LAYER metal3 ;
        RECT 178.800 94.300 179.600 94.400 ;
        RECT 178.800 93.700 197.100 94.300 ;
        RECT 178.800 93.600 179.600 93.700 ;
    END
  END address_b[14]
  PIN address_b[15]
    PORT
      LAYER metal1 ;
        RECT 191.600 111.800 192.400 119.800 ;
        RECT 191.800 109.600 192.400 111.800 ;
        RECT 191.600 102.200 192.400 109.600 ;
      LAYER via1 ;
        RECT 191.600 107.600 192.400 108.400 ;
      LAYER metal2 ;
        RECT 191.600 109.600 192.400 110.400 ;
        RECT 191.700 108.400 192.300 109.600 ;
        RECT 191.600 107.600 192.400 108.400 ;
      LAYER metal3 ;
        RECT 191.600 110.300 192.400 110.400 ;
        RECT 191.600 109.700 197.100 110.300 ;
        RECT 191.600 109.600 192.400 109.700 ;
    END
  END address_b[15]
  OBS
      LAYER metal1 ;
        RECT 2.800 175.200 3.600 179.800 ;
        RECT 6.000 175.200 6.800 179.800 ;
        RECT 9.200 175.200 10.000 179.800 ;
        RECT 12.400 175.200 13.200 179.800 ;
        RECT 15.600 175.400 16.400 179.800 ;
        RECT 19.800 178.400 21.000 179.800 ;
        RECT 19.800 177.800 21.200 178.400 ;
        RECT 24.400 177.800 25.200 179.800 ;
        RECT 28.800 178.400 29.600 179.800 ;
        RECT 28.800 177.800 30.800 178.400 ;
        RECT 20.400 177.000 21.200 177.800 ;
        RECT 24.600 177.200 25.200 177.800 ;
        RECT 24.600 176.600 27.400 177.200 ;
        RECT 26.600 176.400 27.400 176.600 ;
        RECT 28.400 176.400 29.200 177.200 ;
        RECT 30.000 177.000 30.800 177.800 ;
        RECT 18.600 175.400 19.400 175.600 ;
        RECT 2.800 174.400 4.600 175.200 ;
        RECT 6.000 174.400 8.200 175.200 ;
        RECT 9.200 174.400 11.400 175.200 ;
        RECT 12.400 174.400 14.800 175.200 ;
        RECT 3.800 173.800 4.600 174.400 ;
        RECT 7.400 173.800 8.200 174.400 ;
        RECT 10.600 173.800 11.400 174.400 ;
        RECT 3.800 173.000 6.400 173.800 ;
        RECT 7.400 173.000 9.800 173.800 ;
        RECT 10.600 173.000 13.200 173.800 ;
        RECT 3.800 171.600 4.600 173.000 ;
        RECT 7.400 171.600 8.200 173.000 ;
        RECT 10.600 171.600 11.400 173.000 ;
        RECT 14.000 171.600 14.800 174.400 ;
        RECT 2.800 170.800 4.600 171.600 ;
        RECT 6.000 170.800 8.200 171.600 ;
        RECT 9.200 170.800 11.400 171.600 ;
        RECT 12.400 170.800 14.800 171.600 ;
        RECT 15.600 174.800 19.400 175.400 ;
        RECT 15.600 171.400 16.400 174.800 ;
        RECT 22.600 174.200 23.400 174.400 ;
        RECT 26.800 174.200 27.600 174.400 ;
        RECT 28.400 174.200 29.000 176.400 ;
        RECT 33.200 175.000 34.000 179.800 ;
        RECT 34.800 175.200 35.600 179.800 ;
        RECT 34.800 174.600 37.000 175.200 ;
        RECT 39.600 175.000 40.400 179.800 ;
        RECT 44.000 178.400 44.800 179.800 ;
        RECT 42.800 177.800 44.800 178.400 ;
        RECT 48.400 177.800 49.200 179.800 ;
        RECT 52.600 178.400 53.800 179.800 ;
        RECT 52.400 177.800 53.800 178.400 ;
        RECT 42.800 177.000 43.600 177.800 ;
        RECT 48.400 177.200 49.000 177.800 ;
        RECT 44.400 176.400 45.200 177.200 ;
        RECT 46.200 176.600 49.000 177.200 ;
        RECT 52.400 177.000 53.200 177.800 ;
        RECT 46.200 176.400 47.000 176.600 ;
        RECT 31.600 174.200 33.200 174.400 ;
        RECT 22.200 173.600 33.200 174.200 ;
        RECT 20.400 172.800 21.200 173.000 ;
        RECT 17.400 172.200 21.200 172.800 ;
        RECT 17.400 172.000 18.200 172.200 ;
        RECT 19.000 171.400 19.800 171.600 ;
        RECT 15.600 170.800 19.800 171.400 ;
        RECT 2.800 162.200 3.600 170.800 ;
        RECT 6.000 162.200 6.800 170.800 ;
        RECT 9.200 162.200 10.000 170.800 ;
        RECT 12.400 162.200 13.200 170.800 ;
        RECT 15.600 162.200 16.400 170.800 ;
        RECT 22.200 170.400 22.800 173.600 ;
        RECT 29.400 173.400 30.200 173.600 ;
        RECT 28.400 172.400 29.200 172.600 ;
        RECT 31.000 172.400 31.800 172.600 ;
        RECT 26.800 171.800 31.800 172.400 ;
        RECT 26.800 171.600 27.600 171.800 ;
        RECT 34.800 171.600 35.600 173.200 ;
        RECT 36.400 171.600 37.000 174.600 ;
        RECT 40.400 174.200 42.000 174.400 ;
        RECT 44.600 174.200 45.200 176.400 ;
        RECT 54.200 175.400 55.000 175.600 ;
        RECT 57.200 175.400 58.000 179.800 ;
        RECT 54.200 174.800 58.000 175.400 ;
        RECT 50.200 174.200 51.000 174.400 ;
        RECT 40.400 173.600 51.400 174.200 ;
        RECT 43.400 173.400 44.200 173.600 ;
        RECT 41.800 172.400 42.600 172.600 ;
        RECT 41.800 171.800 46.800 172.400 ;
        RECT 46.000 171.600 46.800 171.800 ;
        RECT 28.400 171.000 34.000 171.200 ;
        RECT 28.200 170.800 34.000 171.000 ;
        RECT 20.400 169.800 22.800 170.400 ;
        RECT 24.200 170.600 34.000 170.800 ;
        RECT 24.200 170.200 29.000 170.600 ;
        RECT 20.400 168.800 21.000 169.800 ;
        RECT 19.600 168.000 21.000 168.800 ;
        RECT 22.600 169.000 23.400 169.200 ;
        RECT 24.200 169.000 24.800 170.200 ;
        RECT 22.600 168.400 24.800 169.000 ;
        RECT 25.400 169.000 30.800 169.600 ;
        RECT 25.400 168.800 26.200 169.000 ;
        RECT 30.000 168.800 30.800 169.000 ;
        RECT 23.800 167.400 24.600 167.600 ;
        RECT 26.600 167.400 27.400 167.600 ;
        RECT 20.400 166.200 21.200 167.000 ;
        RECT 23.800 166.800 27.400 167.400 ;
        RECT 24.600 166.200 25.200 166.800 ;
        RECT 30.000 166.200 30.800 167.000 ;
        RECT 19.800 162.200 21.000 166.200 ;
        RECT 24.400 162.200 25.200 166.200 ;
        RECT 28.800 165.600 30.800 166.200 ;
        RECT 28.800 162.200 29.600 165.600 ;
        RECT 33.200 162.200 34.000 170.600 ;
        RECT 36.400 170.800 37.600 171.600 ;
        RECT 39.600 171.000 45.200 171.200 ;
        RECT 39.600 170.800 45.400 171.000 ;
        RECT 36.400 170.200 37.000 170.800 ;
        RECT 34.800 169.600 37.000 170.200 ;
        RECT 39.600 170.600 49.400 170.800 ;
        RECT 34.800 162.200 35.600 169.600 ;
        RECT 39.600 162.200 40.400 170.600 ;
        RECT 44.600 170.200 49.400 170.600 ;
        RECT 42.800 169.000 48.200 169.600 ;
        RECT 42.800 168.800 43.600 169.000 ;
        RECT 47.400 168.800 48.200 169.000 ;
        RECT 48.800 169.000 49.400 170.200 ;
        RECT 50.800 170.400 51.400 173.600 ;
        RECT 52.400 172.800 53.200 173.000 ;
        RECT 52.400 172.200 56.200 172.800 ;
        RECT 55.400 172.000 56.200 172.200 ;
        RECT 53.800 171.400 54.600 171.600 ;
        RECT 57.200 171.400 58.000 174.800 ;
        RECT 63.600 175.200 64.400 179.800 ;
        RECT 68.400 175.200 69.200 179.800 ;
        RECT 73.200 175.200 74.000 179.800 ;
        RECT 78.000 175.400 78.800 179.800 ;
        RECT 82.200 178.400 83.400 179.800 ;
        RECT 82.200 177.800 83.600 178.400 ;
        RECT 86.800 177.800 87.600 179.800 ;
        RECT 91.200 178.400 92.000 179.800 ;
        RECT 91.200 177.800 93.200 178.400 ;
        RECT 82.800 177.000 83.600 177.800 ;
        RECT 87.000 177.200 87.600 177.800 ;
        RECT 87.000 176.600 89.800 177.200 ;
        RECT 89.000 176.400 89.800 176.600 ;
        RECT 90.800 176.400 91.600 177.200 ;
        RECT 92.400 177.000 93.200 177.800 ;
        RECT 81.000 175.400 81.800 175.600 ;
        RECT 63.600 174.600 65.800 175.200 ;
        RECT 68.400 174.600 70.600 175.200 ;
        RECT 73.200 174.600 75.400 175.200 ;
        RECT 63.600 171.600 64.400 173.200 ;
        RECT 65.200 171.600 65.800 174.600 ;
        RECT 68.400 171.600 69.200 173.200 ;
        RECT 70.000 171.600 70.600 174.600 ;
        RECT 73.200 171.600 74.000 173.200 ;
        RECT 74.800 171.600 75.400 174.600 ;
        RECT 78.000 174.800 81.800 175.400 ;
        RECT 53.800 170.800 58.000 171.400 ;
        RECT 50.800 169.800 53.200 170.400 ;
        RECT 50.200 169.000 51.000 169.200 ;
        RECT 48.800 168.400 51.000 169.000 ;
        RECT 52.600 168.800 53.200 169.800 ;
        RECT 52.600 168.000 54.000 168.800 ;
        RECT 46.200 167.400 47.000 167.600 ;
        RECT 49.000 167.400 49.800 167.600 ;
        RECT 42.800 166.200 43.600 167.000 ;
        RECT 46.200 166.800 49.800 167.400 ;
        RECT 48.400 166.200 49.000 166.800 ;
        RECT 52.400 166.200 53.200 167.000 ;
        RECT 42.800 165.600 44.800 166.200 ;
        RECT 44.000 162.200 44.800 165.600 ;
        RECT 48.400 162.200 49.200 166.200 ;
        RECT 52.600 162.200 53.800 166.200 ;
        RECT 57.200 164.300 58.000 170.800 ;
        RECT 65.200 170.800 66.400 171.600 ;
        RECT 70.000 170.800 71.200 171.600 ;
        RECT 74.800 170.800 76.000 171.600 ;
        RECT 78.000 171.400 78.800 174.800 ;
        RECT 85.000 174.200 85.800 174.400 ;
        RECT 90.800 174.200 91.400 176.400 ;
        RECT 95.600 175.000 96.400 179.800 ;
        RECT 100.400 175.200 101.200 179.800 ;
        RECT 105.200 175.200 106.000 179.800 ;
        RECT 99.000 174.600 101.200 175.200 ;
        RECT 103.800 174.600 106.000 175.200 ;
        RECT 106.800 175.400 107.600 179.800 ;
        RECT 111.000 178.400 112.200 179.800 ;
        RECT 111.000 177.800 112.400 178.400 ;
        RECT 115.600 177.800 116.400 179.800 ;
        RECT 120.000 178.400 120.800 179.800 ;
        RECT 120.000 177.800 122.000 178.400 ;
        RECT 111.600 177.000 112.400 177.800 ;
        RECT 115.800 177.200 116.400 177.800 ;
        RECT 115.800 176.600 118.600 177.200 ;
        RECT 117.800 176.400 118.600 176.600 ;
        RECT 119.600 176.400 120.400 177.200 ;
        RECT 121.200 177.000 122.000 177.800 ;
        RECT 109.800 175.400 110.600 175.600 ;
        RECT 106.800 174.800 110.600 175.400 ;
        RECT 94.000 174.200 95.600 174.400 ;
        RECT 84.600 173.600 95.600 174.200 ;
        RECT 82.800 172.800 83.600 173.000 ;
        RECT 79.800 172.200 83.600 172.800 ;
        RECT 79.800 172.000 80.600 172.200 ;
        RECT 81.400 171.400 82.200 171.600 ;
        RECT 78.000 170.800 82.200 171.400 ;
        RECT 65.200 170.200 65.800 170.800 ;
        RECT 70.000 170.200 70.600 170.800 ;
        RECT 74.800 170.200 75.400 170.800 ;
        RECT 63.600 169.600 65.800 170.200 ;
        RECT 68.400 169.600 70.600 170.200 ;
        RECT 73.200 169.600 75.400 170.200 ;
        RECT 58.800 164.300 59.600 164.400 ;
        RECT 57.200 163.700 59.600 164.300 ;
        RECT 57.200 162.200 58.000 163.700 ;
        RECT 58.800 163.600 59.600 163.700 ;
        RECT 63.600 162.200 64.400 169.600 ;
        RECT 68.400 162.200 69.200 169.600 ;
        RECT 73.200 162.200 74.000 169.600 ;
        RECT 78.000 162.200 78.800 170.800 ;
        RECT 84.600 170.400 85.200 173.600 ;
        RECT 91.800 173.400 92.600 173.600 ;
        RECT 90.800 172.400 91.600 172.600 ;
        RECT 93.400 172.400 94.200 172.600 ;
        RECT 89.200 171.800 94.200 172.400 ;
        RECT 89.200 171.600 90.000 171.800 ;
        RECT 99.000 171.600 99.600 174.600 ;
        RECT 100.400 171.600 101.200 173.200 ;
        RECT 103.800 171.600 104.400 174.600 ;
        RECT 105.200 171.600 106.000 173.200 ;
        RECT 90.800 171.000 96.400 171.200 ;
        RECT 90.600 170.800 96.400 171.000 ;
        RECT 98.400 170.800 99.600 171.600 ;
        RECT 103.200 170.800 104.400 171.600 ;
        RECT 82.800 169.800 85.200 170.400 ;
        RECT 86.600 170.600 96.400 170.800 ;
        RECT 86.600 170.200 91.400 170.600 ;
        RECT 82.800 168.800 83.400 169.800 ;
        RECT 82.000 168.000 83.400 168.800 ;
        RECT 85.000 169.000 85.800 169.200 ;
        RECT 86.600 169.000 87.200 170.200 ;
        RECT 85.000 168.400 87.200 169.000 ;
        RECT 87.800 169.000 93.200 169.600 ;
        RECT 87.800 168.800 88.600 169.000 ;
        RECT 92.400 168.800 93.200 169.000 ;
        RECT 86.200 167.400 87.000 167.600 ;
        RECT 89.000 167.400 89.800 167.600 ;
        RECT 82.800 166.200 83.600 167.000 ;
        RECT 86.200 166.800 89.800 167.400 ;
        RECT 87.000 166.200 87.600 166.800 ;
        RECT 92.400 166.200 93.200 167.000 ;
        RECT 82.200 162.200 83.400 166.200 ;
        RECT 86.800 162.200 87.600 166.200 ;
        RECT 91.200 165.600 93.200 166.200 ;
        RECT 91.200 162.200 92.000 165.600 ;
        RECT 95.600 162.200 96.400 170.600 ;
        RECT 99.000 170.200 99.600 170.800 ;
        RECT 103.800 170.200 104.400 170.800 ;
        RECT 106.800 171.400 107.600 174.800 ;
        RECT 113.800 174.200 114.600 174.400 ;
        RECT 119.600 174.200 120.200 176.400 ;
        RECT 124.400 175.000 125.200 179.800 ;
        RECT 126.000 175.200 126.800 179.800 ;
        RECT 130.800 175.200 131.600 179.800 ;
        RECT 140.400 175.400 141.200 179.800 ;
        RECT 144.600 178.400 145.800 179.800 ;
        RECT 144.600 177.800 146.000 178.400 ;
        RECT 149.200 177.800 150.000 179.800 ;
        RECT 153.600 178.400 154.400 179.800 ;
        RECT 153.600 177.800 155.600 178.400 ;
        RECT 145.200 177.000 146.000 177.800 ;
        RECT 149.400 177.200 150.000 177.800 ;
        RECT 149.400 176.600 152.200 177.200 ;
        RECT 151.400 176.400 152.200 176.600 ;
        RECT 153.200 176.400 154.000 177.200 ;
        RECT 154.800 177.000 155.600 177.800 ;
        RECT 143.400 175.400 144.200 175.600 ;
        RECT 126.000 174.600 128.200 175.200 ;
        RECT 130.800 174.600 133.000 175.200 ;
        RECT 122.800 174.200 124.400 174.400 ;
        RECT 113.400 173.600 124.400 174.200 ;
        RECT 111.600 172.800 112.400 173.000 ;
        RECT 108.600 172.200 112.400 172.800 ;
        RECT 113.400 172.400 114.000 173.600 ;
        RECT 120.600 173.400 121.400 173.600 ;
        RECT 119.600 172.400 120.400 172.600 ;
        RECT 122.200 172.400 123.000 172.600 ;
        RECT 108.600 172.000 109.400 172.200 ;
        RECT 113.200 171.600 114.000 172.400 ;
        RECT 118.000 171.800 123.000 172.400 ;
        RECT 118.000 171.600 118.800 171.800 ;
        RECT 126.000 171.600 126.800 173.200 ;
        RECT 127.600 171.600 128.200 174.600 ;
        RECT 130.800 171.600 131.600 173.200 ;
        RECT 132.400 171.600 133.000 174.600 ;
        RECT 140.400 174.800 144.200 175.400 ;
        RECT 110.200 171.400 111.000 171.600 ;
        RECT 106.800 170.800 111.000 171.400 ;
        RECT 99.000 169.600 101.200 170.200 ;
        RECT 103.800 169.600 106.000 170.200 ;
        RECT 100.400 162.200 101.200 169.600 ;
        RECT 105.200 162.200 106.000 169.600 ;
        RECT 106.800 162.200 107.600 170.800 ;
        RECT 113.400 170.400 114.000 171.600 ;
        RECT 119.600 171.000 125.200 171.200 ;
        RECT 119.400 170.800 125.200 171.000 ;
        RECT 111.600 169.800 114.000 170.400 ;
        RECT 115.400 170.600 125.200 170.800 ;
        RECT 115.400 170.200 120.200 170.600 ;
        RECT 111.600 168.800 112.200 169.800 ;
        RECT 110.800 168.000 112.200 168.800 ;
        RECT 113.800 169.000 114.600 169.200 ;
        RECT 115.400 169.000 116.000 170.200 ;
        RECT 113.800 168.400 116.000 169.000 ;
        RECT 116.600 169.000 122.000 169.600 ;
        RECT 116.600 168.800 117.400 169.000 ;
        RECT 121.200 168.800 122.000 169.000 ;
        RECT 115.000 167.400 115.800 167.600 ;
        RECT 117.800 167.400 118.600 167.600 ;
        RECT 111.600 166.200 112.400 167.000 ;
        RECT 115.000 166.800 118.600 167.400 ;
        RECT 115.800 166.200 116.400 166.800 ;
        RECT 121.200 166.200 122.000 167.000 ;
        RECT 111.000 162.200 112.200 166.200 ;
        RECT 115.600 162.200 116.400 166.200 ;
        RECT 120.000 165.600 122.000 166.200 ;
        RECT 120.000 162.200 120.800 165.600 ;
        RECT 124.400 162.200 125.200 170.600 ;
        RECT 127.600 170.800 128.800 171.600 ;
        RECT 132.400 170.800 133.600 171.600 ;
        RECT 140.400 171.400 141.200 174.800 ;
        RECT 147.400 174.200 148.200 174.400 ;
        RECT 153.200 174.200 153.800 176.400 ;
        RECT 158.000 175.000 158.800 179.800 ;
        RECT 159.600 175.200 160.400 179.800 ;
        RECT 159.600 174.600 161.800 175.200 ;
        RECT 164.400 175.000 165.200 179.800 ;
        RECT 168.800 178.400 169.600 179.800 ;
        RECT 167.600 177.800 169.600 178.400 ;
        RECT 173.200 177.800 174.000 179.800 ;
        RECT 177.400 178.400 178.600 179.800 ;
        RECT 177.200 177.800 178.600 178.400 ;
        RECT 167.600 177.000 168.400 177.800 ;
        RECT 173.200 177.200 173.800 177.800 ;
        RECT 169.200 176.400 170.000 177.200 ;
        RECT 171.000 176.600 173.800 177.200 ;
        RECT 177.200 177.000 178.000 177.800 ;
        RECT 171.000 176.400 171.800 176.600 ;
        RECT 156.400 174.200 158.000 174.400 ;
        RECT 147.000 173.600 158.000 174.200 ;
        RECT 145.200 172.800 146.000 173.000 ;
        RECT 142.200 172.200 146.000 172.800 ;
        RECT 147.000 172.400 147.600 173.600 ;
        RECT 154.200 173.400 155.000 173.600 ;
        RECT 153.200 172.400 154.000 172.600 ;
        RECT 155.800 172.400 156.600 172.600 ;
        RECT 142.200 172.000 143.000 172.200 ;
        RECT 146.800 171.600 147.600 172.400 ;
        RECT 151.600 171.800 156.600 172.400 ;
        RECT 151.600 171.600 152.400 171.800 ;
        RECT 159.600 171.600 160.400 173.200 ;
        RECT 161.200 171.600 161.800 174.600 ;
        RECT 165.200 174.200 166.800 174.400 ;
        RECT 169.400 174.200 170.000 176.400 ;
        RECT 179.000 175.400 179.800 175.600 ;
        RECT 182.000 175.400 182.800 179.800 ;
        RECT 179.000 174.800 182.800 175.400 ;
        RECT 175.000 174.200 175.800 174.400 ;
        RECT 165.200 173.600 176.200 174.200 ;
        RECT 168.200 173.400 169.000 173.600 ;
        RECT 166.600 172.400 167.400 172.600 ;
        RECT 166.600 171.800 171.600 172.400 ;
        RECT 170.800 171.600 171.600 171.800 ;
        RECT 143.800 171.400 144.600 171.600 ;
        RECT 140.400 170.800 144.600 171.400 ;
        RECT 127.600 170.200 128.200 170.800 ;
        RECT 132.400 170.200 133.000 170.800 ;
        RECT 126.000 169.600 128.200 170.200 ;
        RECT 130.800 169.600 133.000 170.200 ;
        RECT 126.000 162.200 126.800 169.600 ;
        RECT 130.800 162.200 131.600 169.600 ;
        RECT 140.400 162.200 141.200 170.800 ;
        RECT 147.000 170.400 147.600 171.600 ;
        RECT 153.200 171.000 158.800 171.200 ;
        RECT 153.000 170.800 158.800 171.000 ;
        RECT 145.200 169.800 147.600 170.400 ;
        RECT 149.000 170.600 158.800 170.800 ;
        RECT 149.000 170.200 153.800 170.600 ;
        RECT 145.200 168.800 145.800 169.800 ;
        RECT 144.400 168.000 145.800 168.800 ;
        RECT 147.400 169.000 148.200 169.200 ;
        RECT 149.000 169.000 149.600 170.200 ;
        RECT 147.400 168.400 149.600 169.000 ;
        RECT 150.200 169.000 155.600 169.600 ;
        RECT 150.200 168.800 151.000 169.000 ;
        RECT 154.800 168.800 155.600 169.000 ;
        RECT 148.600 167.400 149.400 167.600 ;
        RECT 151.400 167.400 152.200 167.600 ;
        RECT 145.200 166.200 146.000 167.000 ;
        RECT 148.600 166.800 152.200 167.400 ;
        RECT 149.400 166.200 150.000 166.800 ;
        RECT 154.800 166.200 155.600 167.000 ;
        RECT 144.600 162.200 145.800 166.200 ;
        RECT 149.200 162.200 150.000 166.200 ;
        RECT 153.600 165.600 155.600 166.200 ;
        RECT 153.600 162.200 154.400 165.600 ;
        RECT 158.000 162.200 158.800 170.600 ;
        RECT 161.200 170.800 162.400 171.600 ;
        RECT 164.400 171.000 170.000 171.200 ;
        RECT 164.400 170.800 170.200 171.000 ;
        RECT 161.200 170.200 161.800 170.800 ;
        RECT 159.600 169.600 161.800 170.200 ;
        RECT 164.400 170.600 174.200 170.800 ;
        RECT 159.600 162.200 160.400 169.600 ;
        RECT 164.400 162.200 165.200 170.600 ;
        RECT 169.400 170.200 174.200 170.600 ;
        RECT 167.600 169.000 173.000 169.600 ;
        RECT 167.600 168.800 168.400 169.000 ;
        RECT 172.200 168.800 173.000 169.000 ;
        RECT 173.600 169.000 174.200 170.200 ;
        RECT 175.600 170.400 176.200 173.600 ;
        RECT 177.200 172.800 178.000 173.000 ;
        RECT 177.200 172.200 181.000 172.800 ;
        RECT 180.200 172.000 181.000 172.200 ;
        RECT 178.600 171.400 179.400 171.600 ;
        RECT 182.000 171.400 182.800 174.800 ;
        RECT 178.600 170.800 182.800 171.400 ;
        RECT 175.600 169.800 178.000 170.400 ;
        RECT 175.000 169.000 175.800 169.200 ;
        RECT 173.600 168.400 175.800 169.000 ;
        RECT 177.400 168.800 178.000 169.800 ;
        RECT 177.400 168.000 178.800 168.800 ;
        RECT 171.000 167.400 171.800 167.600 ;
        RECT 173.800 167.400 174.600 167.600 ;
        RECT 167.600 166.200 168.400 167.000 ;
        RECT 171.000 166.800 174.600 167.400 ;
        RECT 173.200 166.200 173.800 166.800 ;
        RECT 177.200 166.200 178.000 167.000 ;
        RECT 167.600 165.600 169.600 166.200 ;
        RECT 168.800 162.200 169.600 165.600 ;
        RECT 173.200 162.200 174.000 166.200 ;
        RECT 177.400 162.200 178.600 166.200 ;
        RECT 182.000 162.200 182.800 170.800 ;
        RECT 183.600 175.800 184.400 179.800 ;
        RECT 186.800 177.800 187.600 179.800 ;
        RECT 183.600 172.400 184.200 175.800 ;
        RECT 186.800 175.600 187.400 177.800 ;
        RECT 185.000 175.000 187.400 175.600 ;
        RECT 190.000 175.200 190.800 179.800 ;
        RECT 183.600 171.600 184.400 172.400 ;
        RECT 185.000 172.000 185.600 175.000 ;
        RECT 190.000 174.600 192.200 175.200 ;
        RECT 186.600 174.300 187.600 174.400 ;
        RECT 188.400 174.300 189.200 174.400 ;
        RECT 186.600 173.700 189.200 174.300 ;
        RECT 186.600 173.600 187.600 173.700 ;
        RECT 188.400 173.600 189.200 173.700 ;
        RECT 186.400 172.800 187.200 173.600 ;
        RECT 183.600 170.200 184.200 171.600 ;
        RECT 185.000 171.400 185.800 172.000 ;
        RECT 190.000 171.600 190.800 173.200 ;
        RECT 191.600 171.600 192.200 174.600 ;
        RECT 185.000 171.200 189.200 171.400 ;
        RECT 185.200 170.800 189.200 171.200 ;
        RECT 183.600 169.600 185.000 170.200 ;
        RECT 184.200 162.200 185.000 169.600 ;
        RECT 188.400 162.200 189.200 170.800 ;
        RECT 191.600 170.800 192.800 171.600 ;
        RECT 191.600 170.200 192.200 170.800 ;
        RECT 190.000 169.600 192.200 170.200 ;
        RECT 190.000 162.200 190.800 169.600 ;
        RECT 1.200 151.200 2.000 159.800 ;
        RECT 5.400 155.800 6.600 159.800 ;
        RECT 10.000 155.800 10.800 159.800 ;
        RECT 14.400 156.400 15.200 159.800 ;
        RECT 14.400 155.800 16.400 156.400 ;
        RECT 6.000 155.000 6.800 155.800 ;
        RECT 10.200 155.200 10.800 155.800 ;
        RECT 9.400 154.600 13.000 155.200 ;
        RECT 15.600 155.000 16.400 155.800 ;
        RECT 9.400 154.400 10.200 154.600 ;
        RECT 12.200 154.400 13.000 154.600 ;
        RECT 5.200 153.200 6.600 154.000 ;
        RECT 6.000 152.200 6.600 153.200 ;
        RECT 8.200 153.000 10.400 153.600 ;
        RECT 8.200 152.800 9.000 153.000 ;
        RECT 6.000 151.600 8.400 152.200 ;
        RECT 1.200 150.600 5.400 151.200 ;
        RECT 1.200 147.200 2.000 150.600 ;
        RECT 4.600 150.400 5.400 150.600 ;
        RECT 3.000 149.800 3.800 150.000 ;
        RECT 3.000 149.200 6.800 149.800 ;
        RECT 6.000 149.000 6.800 149.200 ;
        RECT 7.800 148.400 8.400 151.600 ;
        RECT 9.800 151.800 10.400 153.000 ;
        RECT 11.000 153.000 11.800 153.200 ;
        RECT 15.600 153.000 16.400 153.200 ;
        RECT 11.000 152.400 16.400 153.000 ;
        RECT 9.800 151.400 14.600 151.800 ;
        RECT 18.800 151.400 19.600 159.800 ;
        RECT 9.800 151.200 19.600 151.400 ;
        RECT 13.800 151.000 19.600 151.200 ;
        RECT 14.000 150.800 19.600 151.000 ;
        RECT 20.400 151.200 21.200 159.800 ;
        RECT 24.600 155.800 25.800 159.800 ;
        RECT 29.200 155.800 30.000 159.800 ;
        RECT 33.600 156.400 34.400 159.800 ;
        RECT 33.600 155.800 35.600 156.400 ;
        RECT 25.200 155.000 26.000 155.800 ;
        RECT 29.400 155.200 30.000 155.800 ;
        RECT 28.600 154.600 32.200 155.200 ;
        RECT 34.800 155.000 35.600 155.800 ;
        RECT 28.600 154.400 29.400 154.600 ;
        RECT 31.400 154.400 32.200 154.600 ;
        RECT 24.400 153.200 25.800 154.000 ;
        RECT 25.200 152.200 25.800 153.200 ;
        RECT 27.400 153.000 29.600 153.600 ;
        RECT 27.400 152.800 28.200 153.000 ;
        RECT 25.200 151.600 27.600 152.200 ;
        RECT 20.400 150.600 24.600 151.200 ;
        RECT 12.400 150.200 13.200 150.400 ;
        RECT 12.400 149.600 17.400 150.200 ;
        RECT 14.000 149.400 14.800 149.600 ;
        RECT 16.600 149.400 17.400 149.600 ;
        RECT 15.000 148.400 15.800 148.600 ;
        RECT 7.800 147.800 18.800 148.400 ;
        RECT 8.200 147.600 9.000 147.800 ;
        RECT 12.400 147.600 13.200 147.800 ;
        RECT 1.200 146.600 5.000 147.200 ;
        RECT 1.200 142.200 2.000 146.600 ;
        RECT 4.200 146.400 5.000 146.600 ;
        RECT 14.000 145.600 14.600 147.800 ;
        RECT 17.200 147.600 18.800 147.800 ;
        RECT 20.400 147.200 21.200 150.600 ;
        RECT 23.800 150.400 24.600 150.600 ;
        RECT 27.000 150.400 27.600 151.600 ;
        RECT 29.000 151.800 29.600 153.000 ;
        RECT 30.200 153.000 31.000 153.200 ;
        RECT 34.800 153.000 35.600 153.200 ;
        RECT 30.200 152.400 35.600 153.000 ;
        RECT 29.000 151.400 33.800 151.800 ;
        RECT 38.000 151.400 38.800 159.800 ;
        RECT 29.000 151.200 38.800 151.400 ;
        RECT 33.000 151.000 38.800 151.200 ;
        RECT 33.200 150.800 38.800 151.000 ;
        RECT 39.600 151.800 40.400 159.800 ;
        RECT 42.800 155.800 43.600 159.800 ;
        RECT 39.600 150.400 40.200 151.800 ;
        RECT 42.800 151.600 43.400 155.800 ;
        RECT 41.000 151.000 43.400 151.600 ;
        RECT 22.200 149.800 23.000 150.000 ;
        RECT 22.200 149.200 26.000 149.800 ;
        RECT 26.800 149.600 27.600 150.400 ;
        RECT 31.600 150.200 32.400 150.400 ;
        RECT 31.600 149.600 36.600 150.200 ;
        RECT 25.200 149.000 26.000 149.200 ;
        RECT 27.000 148.400 27.600 149.600 ;
        RECT 33.200 149.400 34.000 149.600 ;
        RECT 35.800 149.400 36.600 149.600 ;
        RECT 39.600 149.600 40.400 150.400 ;
        RECT 34.200 148.400 35.000 148.600 ;
        RECT 27.000 147.800 38.000 148.400 ;
        RECT 27.400 147.600 28.200 147.800 ;
        RECT 12.200 145.400 13.000 145.600 ;
        RECT 6.000 144.200 6.800 145.000 ;
        RECT 10.200 144.800 13.000 145.400 ;
        RECT 14.000 144.800 14.800 145.600 ;
        RECT 10.200 144.200 10.800 144.800 ;
        RECT 15.600 144.200 16.400 145.000 ;
        RECT 5.400 143.600 6.800 144.200 ;
        RECT 5.400 142.200 6.600 143.600 ;
        RECT 10.000 142.200 10.800 144.200 ;
        RECT 14.400 143.600 16.400 144.200 ;
        RECT 14.400 142.200 15.200 143.600 ;
        RECT 18.800 142.200 19.600 147.000 ;
        RECT 20.400 146.600 24.200 147.200 ;
        RECT 20.400 142.200 21.200 146.600 ;
        RECT 23.400 146.400 24.200 146.600 ;
        RECT 33.200 145.600 33.800 147.800 ;
        RECT 36.400 147.600 38.000 147.800 ;
        RECT 31.400 145.400 32.200 145.600 ;
        RECT 25.200 144.200 26.000 145.000 ;
        RECT 29.400 144.800 32.200 145.400 ;
        RECT 33.200 144.800 34.000 145.600 ;
        RECT 29.400 144.200 30.000 144.800 ;
        RECT 34.800 144.200 35.600 145.000 ;
        RECT 24.600 143.600 26.000 144.200 ;
        RECT 24.600 142.200 25.800 143.600 ;
        RECT 29.200 142.200 30.000 144.200 ;
        RECT 33.600 143.600 35.600 144.200 ;
        RECT 33.600 142.200 34.400 143.600 ;
        RECT 38.000 142.200 38.800 147.000 ;
        RECT 39.600 146.200 40.200 149.600 ;
        RECT 41.000 147.600 41.600 151.000 ;
        RECT 42.800 149.600 43.600 150.400 ;
        RECT 42.800 148.800 43.400 149.600 ;
        RECT 42.400 148.000 43.600 148.800 ;
        RECT 44.400 147.600 45.200 149.200 ;
        RECT 47.600 148.300 48.400 159.800 ;
        RECT 49.200 152.400 50.000 159.800 ;
        RECT 52.400 152.400 53.200 159.800 ;
        RECT 49.200 151.800 53.200 152.400 ;
        RECT 54.000 151.800 54.800 159.800 ;
        RECT 50.000 150.400 50.800 150.800 ;
        RECT 54.000 150.400 54.600 151.800 ;
        RECT 49.200 149.800 50.800 150.400 ;
        RECT 52.400 149.800 54.800 150.400 ;
        RECT 49.200 149.600 50.000 149.800 ;
        RECT 52.400 149.600 53.200 149.800 ;
        RECT 54.000 149.600 54.800 149.800 ;
        RECT 50.800 148.300 51.600 149.200 ;
        RECT 47.600 147.700 51.600 148.300 ;
        RECT 40.800 147.400 41.600 147.600 ;
        RECT 40.800 147.000 43.800 147.400 ;
        RECT 40.800 146.800 45.000 147.000 ;
        RECT 43.200 146.400 45.000 146.800 ;
        RECT 44.400 146.200 45.000 146.400 ;
        RECT 39.600 145.200 41.000 146.200 ;
        RECT 40.200 142.200 41.000 145.200 ;
        RECT 44.400 142.200 45.200 146.200 ;
        RECT 46.000 144.800 46.800 146.400 ;
        RECT 47.600 142.200 48.400 147.700 ;
        RECT 50.800 147.600 51.600 147.700 ;
        RECT 52.400 146.200 53.000 149.600 ;
        RECT 58.800 148.300 59.600 148.400 ;
        RECT 60.400 148.300 61.200 148.400 ;
        RECT 58.800 147.700 61.200 148.300 ;
        RECT 58.800 147.600 59.600 147.700 ;
        RECT 60.400 146.800 61.200 147.700 ;
        RECT 52.400 142.200 53.200 146.200 ;
        RECT 54.000 145.600 54.800 146.400 ;
        RECT 62.000 146.200 62.800 159.800 ;
        RECT 63.600 151.600 64.400 153.200 ;
        RECT 66.800 148.300 67.600 159.800 ;
        RECT 68.400 151.800 69.200 159.800 ;
        RECT 70.000 152.400 70.800 159.800 ;
        RECT 73.200 152.400 74.000 159.800 ;
        RECT 70.000 151.800 74.000 152.400 ;
        RECT 68.600 150.400 69.200 151.800 ;
        RECT 74.800 151.600 75.600 153.200 ;
        RECT 72.400 150.400 73.200 150.800 ;
        RECT 68.400 149.800 70.800 150.400 ;
        RECT 72.400 149.800 74.000 150.400 ;
        RECT 68.400 149.600 69.200 149.800 ;
        RECT 70.000 149.600 70.800 149.800 ;
        RECT 73.200 149.600 74.000 149.800 ;
        RECT 68.400 148.300 69.200 148.400 ;
        RECT 66.800 147.700 69.200 148.300 ;
        RECT 62.000 145.600 63.800 146.200 ;
        RECT 53.800 144.800 54.600 145.600 ;
        RECT 63.000 144.400 63.800 145.600 ;
        RECT 65.200 144.800 66.000 146.400 ;
        RECT 63.000 143.600 64.400 144.400 ;
        RECT 63.000 142.200 63.800 143.600 ;
        RECT 66.800 142.200 67.600 147.700 ;
        RECT 68.400 147.600 69.200 147.700 ;
        RECT 68.400 145.600 69.200 146.400 ;
        RECT 70.200 146.200 70.800 149.600 ;
        RECT 71.600 147.600 72.400 149.200 ;
        RECT 76.400 146.200 77.200 159.800 ;
        RECT 78.000 148.300 78.800 148.400 ;
        RECT 78.000 147.700 80.300 148.300 ;
        RECT 78.000 146.800 78.800 147.700 ;
        RECT 79.700 146.400 80.300 147.700 ;
        RECT 68.600 144.800 69.400 145.600 ;
        RECT 70.000 142.200 70.800 146.200 ;
        RECT 75.400 145.600 77.200 146.200 ;
        RECT 75.400 144.400 76.200 145.600 ;
        RECT 79.600 144.800 80.400 146.400 ;
        RECT 74.800 143.600 76.200 144.400 ;
        RECT 75.400 142.200 76.200 143.600 ;
        RECT 81.200 142.200 82.000 159.800 ;
        RECT 83.400 152.400 84.200 159.800 ;
        RECT 82.800 151.800 84.200 152.400 ;
        RECT 82.800 150.400 83.400 151.800 ;
        RECT 87.600 151.200 88.400 159.800 ;
        RECT 89.200 152.400 90.000 159.800 ;
        RECT 92.400 152.400 93.200 159.800 ;
        RECT 89.200 151.800 93.200 152.400 ;
        RECT 94.000 152.300 94.800 159.800 ;
        RECT 97.200 155.800 98.000 159.800 ;
        RECT 95.600 152.300 96.400 152.400 ;
        RECT 84.400 150.800 88.400 151.200 ;
        RECT 94.000 151.700 96.400 152.300 ;
        RECT 84.200 150.600 88.400 150.800 ;
        RECT 82.800 149.600 83.600 150.400 ;
        RECT 84.200 150.000 85.000 150.600 ;
        RECT 90.000 150.400 90.800 150.800 ;
        RECT 94.000 150.400 94.600 151.700 ;
        RECT 95.600 151.600 96.400 151.700 ;
        RECT 97.400 151.600 98.000 155.800 ;
        RECT 100.400 151.800 101.200 159.800 ;
        RECT 97.400 151.000 99.800 151.600 ;
        RECT 82.800 146.200 83.400 149.600 ;
        RECT 84.200 147.000 84.800 150.000 ;
        RECT 89.200 149.800 90.800 150.400 ;
        RECT 92.400 149.800 94.800 150.400 ;
        RECT 89.200 149.600 90.000 149.800 ;
        RECT 85.600 148.400 86.400 149.200 ;
        RECT 85.800 148.300 86.800 148.400 ;
        RECT 90.800 148.300 91.600 149.200 ;
        RECT 85.800 147.700 91.600 148.300 ;
        RECT 85.800 147.600 86.800 147.700 ;
        RECT 90.800 147.600 91.600 147.700 ;
        RECT 84.200 146.400 86.600 147.000 ;
        RECT 82.800 142.200 83.600 146.200 ;
        RECT 86.000 144.200 86.600 146.400 ;
        RECT 87.600 144.800 88.400 146.400 ;
        RECT 92.400 146.200 93.000 149.800 ;
        RECT 94.000 149.600 94.800 149.800 ;
        RECT 97.200 149.600 98.000 150.400 ;
        RECT 94.000 148.300 94.800 148.400 ;
        RECT 95.600 148.300 96.400 149.200 ;
        RECT 94.000 147.700 96.400 148.300 ;
        RECT 97.400 148.800 98.000 149.600 ;
        RECT 97.400 148.200 98.400 148.800 ;
        RECT 97.600 148.000 98.400 148.200 ;
        RECT 94.000 147.600 94.800 147.700 ;
        RECT 95.600 147.600 96.400 147.700 ;
        RECT 99.200 147.600 99.800 151.000 ;
        RECT 100.600 150.400 101.200 151.800 ;
        RECT 103.600 151.200 104.400 159.800 ;
        RECT 106.800 151.200 107.600 159.800 ;
        RECT 110.000 151.200 110.800 159.800 ;
        RECT 113.200 151.200 114.000 159.800 ;
        RECT 116.400 152.400 117.200 159.800 ;
        RECT 119.600 152.400 120.400 159.800 ;
        RECT 116.400 151.800 120.400 152.400 ;
        RECT 121.200 151.800 122.000 159.800 ;
        RECT 123.600 153.600 124.400 154.400 ;
        RECT 123.600 152.400 124.200 153.600 ;
        RECT 125.000 152.400 125.800 159.800 ;
        RECT 122.800 151.800 124.200 152.400 ;
        RECT 124.800 151.800 125.800 152.400 ;
        RECT 103.600 150.400 105.400 151.200 ;
        RECT 106.800 150.400 109.000 151.200 ;
        RECT 110.000 150.400 112.200 151.200 ;
        RECT 113.200 150.400 115.600 151.200 ;
        RECT 117.200 150.400 118.000 150.800 ;
        RECT 121.200 150.400 121.800 151.800 ;
        RECT 122.800 151.600 123.600 151.800 ;
        RECT 100.400 149.600 101.200 150.400 ;
        RECT 99.200 147.400 100.000 147.600 ;
        RECT 97.000 147.000 100.000 147.400 ;
        RECT 95.800 146.800 100.000 147.000 ;
        RECT 95.800 146.400 97.600 146.800 ;
        RECT 95.800 146.200 96.400 146.400 ;
        RECT 100.600 146.200 101.200 149.600 ;
        RECT 104.600 149.000 105.400 150.400 ;
        RECT 108.200 149.000 109.000 150.400 ;
        RECT 111.400 149.000 112.200 150.400 ;
        RECT 104.600 148.200 107.200 149.000 ;
        RECT 108.200 148.200 110.600 149.000 ;
        RECT 111.400 148.200 114.000 149.000 ;
        RECT 104.600 147.600 105.400 148.200 ;
        RECT 108.200 147.600 109.000 148.200 ;
        RECT 111.400 147.600 112.200 148.200 ;
        RECT 114.800 147.600 115.600 150.400 ;
        RECT 116.400 149.800 118.000 150.400 ;
        RECT 119.600 149.800 122.000 150.400 ;
        RECT 116.400 149.600 117.200 149.800 ;
        RECT 119.600 149.600 120.400 149.800 ;
        RECT 121.200 149.600 122.000 149.800 ;
        RECT 118.000 147.600 118.800 149.200 ;
        RECT 86.000 142.200 86.800 144.200 ;
        RECT 92.400 142.200 93.200 146.200 ;
        RECT 95.600 142.200 96.400 146.200 ;
        RECT 99.800 145.200 101.200 146.200 ;
        RECT 103.600 146.800 105.400 147.600 ;
        RECT 106.800 146.800 109.000 147.600 ;
        RECT 110.000 146.800 112.200 147.600 ;
        RECT 113.200 146.800 115.600 147.600 ;
        RECT 99.800 142.200 100.600 145.200 ;
        RECT 103.600 142.200 104.400 146.800 ;
        RECT 106.800 142.200 107.600 146.800 ;
        RECT 110.000 142.200 110.800 146.800 ;
        RECT 113.200 142.200 114.000 146.800 ;
        RECT 119.600 146.200 120.200 149.600 ;
        RECT 124.800 148.400 125.400 151.800 ;
        RECT 126.000 148.800 126.800 150.400 ;
        RECT 122.800 147.600 125.400 148.400 ;
        RECT 127.600 148.300 128.400 148.400 ;
        RECT 129.200 148.300 130.000 148.400 ;
        RECT 127.600 148.200 130.000 148.300 ;
        RECT 126.800 147.700 130.000 148.200 ;
        RECT 126.800 147.600 128.400 147.700 ;
        RECT 121.200 146.300 122.000 146.400 ;
        RECT 123.000 146.300 123.600 147.600 ;
        RECT 126.800 147.200 127.600 147.600 ;
        RECT 129.200 146.800 130.000 147.700 ;
        RECT 130.800 148.300 131.600 159.800 ;
        RECT 132.400 151.600 133.200 153.200 ;
        RECT 138.800 152.400 139.600 159.800 ;
        RECT 142.000 152.400 142.800 159.800 ;
        RECT 138.800 151.800 142.800 152.400 ;
        RECT 143.600 151.800 144.400 159.800 ;
        RECT 147.800 152.400 148.600 159.800 ;
        RECT 149.200 153.600 150.000 154.400 ;
        RECT 149.400 152.400 150.000 153.600 ;
        RECT 152.200 152.600 153.000 159.800 ;
        RECT 147.800 151.800 148.800 152.400 ;
        RECT 149.400 151.800 150.800 152.400 ;
        RECT 152.200 151.800 154.000 152.600 ;
        RECT 139.600 150.400 140.400 150.800 ;
        RECT 143.600 150.400 144.200 151.800 ;
        RECT 137.200 150.300 138.000 150.400 ;
        RECT 138.800 150.300 140.400 150.400 ;
        RECT 137.200 149.800 140.400 150.300 ;
        RECT 142.000 149.800 144.400 150.400 ;
        RECT 137.200 149.700 139.600 149.800 ;
        RECT 137.200 149.600 138.000 149.700 ;
        RECT 138.800 149.600 139.600 149.700 ;
        RECT 138.800 148.300 139.600 148.400 ;
        RECT 130.800 147.700 139.600 148.300 ;
        RECT 119.600 142.200 120.400 146.200 ;
        RECT 121.200 145.700 123.600 146.300 ;
        RECT 124.600 146.200 128.200 146.600 ;
        RECT 130.800 146.200 131.600 147.700 ;
        RECT 138.800 147.600 139.600 147.700 ;
        RECT 140.400 147.600 141.200 149.200 ;
        RECT 142.000 148.300 142.600 149.800 ;
        RECT 143.600 149.600 144.400 149.800 ;
        RECT 146.800 148.800 147.600 150.400 ;
        RECT 148.200 150.300 148.800 151.800 ;
        RECT 150.000 151.600 150.800 151.800 ;
        RECT 151.600 150.300 152.400 151.200 ;
        RECT 148.200 149.700 152.400 150.300 ;
        RECT 148.200 148.400 148.800 149.700 ;
        RECT 151.600 149.600 152.400 149.700 ;
        RECT 153.200 150.300 153.800 151.800 ;
        RECT 156.400 151.200 157.200 159.800 ;
        RECT 160.600 155.800 161.800 159.800 ;
        RECT 165.200 155.800 166.000 159.800 ;
        RECT 169.600 156.400 170.400 159.800 ;
        RECT 169.600 155.800 171.600 156.400 ;
        RECT 161.200 155.000 162.000 155.800 ;
        RECT 165.400 155.200 166.000 155.800 ;
        RECT 164.600 154.600 168.200 155.200 ;
        RECT 170.800 155.000 171.600 155.800 ;
        RECT 164.600 154.400 165.400 154.600 ;
        RECT 167.400 154.400 168.200 154.600 ;
        RECT 160.400 153.200 161.800 154.000 ;
        RECT 159.600 151.200 160.400 152.400 ;
        RECT 161.200 152.200 161.800 153.200 ;
        RECT 163.400 153.000 165.600 153.600 ;
        RECT 163.400 152.800 164.200 153.000 ;
        RECT 161.200 151.600 163.600 152.200 ;
        RECT 156.400 150.600 160.600 151.200 ;
        RECT 154.800 150.300 155.600 150.400 ;
        RECT 153.200 149.700 155.600 150.300 ;
        RECT 153.200 148.400 153.800 149.700 ;
        RECT 154.800 149.600 155.600 149.700 ;
        RECT 143.600 148.300 144.400 148.400 ;
        RECT 142.000 147.700 144.400 148.300 ;
        RECT 142.000 146.200 142.600 147.700 ;
        RECT 143.600 147.600 144.400 147.700 ;
        RECT 145.200 148.200 146.000 148.400 ;
        RECT 145.200 147.600 146.800 148.200 ;
        RECT 148.200 147.600 150.800 148.400 ;
        RECT 153.200 147.600 154.000 148.400 ;
        RECT 146.000 147.200 146.800 147.600 ;
        RECT 121.200 145.600 122.000 145.700 ;
        RECT 121.000 144.800 121.800 145.600 ;
        RECT 122.800 142.200 123.600 145.700 ;
        RECT 124.400 146.000 128.400 146.200 ;
        RECT 124.400 142.200 125.200 146.000 ;
        RECT 127.600 142.200 128.400 146.000 ;
        RECT 130.800 145.600 132.600 146.200 ;
        RECT 131.800 142.200 132.600 145.600 ;
        RECT 142.000 142.200 142.800 146.200 ;
        RECT 143.600 145.600 144.400 146.400 ;
        RECT 145.400 146.200 149.000 146.600 ;
        RECT 150.000 146.200 150.600 147.600 ;
        RECT 145.200 146.000 149.200 146.200 ;
        RECT 143.400 144.800 144.200 145.600 ;
        RECT 145.200 142.200 146.000 146.000 ;
        RECT 148.400 142.200 149.200 146.000 ;
        RECT 150.000 142.200 150.800 146.200 ;
        RECT 153.200 144.200 153.800 147.600 ;
        RECT 156.400 147.200 157.200 150.600 ;
        RECT 159.800 150.400 160.600 150.600 ;
        RECT 163.000 150.400 163.600 151.600 ;
        RECT 165.000 151.800 165.600 153.000 ;
        RECT 166.200 153.000 167.000 153.200 ;
        RECT 170.800 153.000 171.600 153.200 ;
        RECT 166.200 152.400 171.600 153.000 ;
        RECT 165.000 151.400 169.800 151.800 ;
        RECT 174.000 151.400 174.800 159.800 ;
        RECT 165.000 151.200 174.800 151.400 ;
        RECT 169.000 151.000 174.800 151.200 ;
        RECT 169.200 150.800 174.800 151.000 ;
        RECT 175.600 151.400 176.400 159.800 ;
        RECT 180.000 156.400 180.800 159.800 ;
        RECT 178.800 155.800 180.800 156.400 ;
        RECT 184.400 155.800 185.200 159.800 ;
        RECT 188.600 155.800 189.800 159.800 ;
        RECT 178.800 155.000 179.600 155.800 ;
        RECT 184.400 155.200 185.000 155.800 ;
        RECT 182.200 154.600 185.800 155.200 ;
        RECT 188.400 155.000 189.200 155.800 ;
        RECT 182.200 154.400 183.000 154.600 ;
        RECT 185.000 154.400 185.800 154.600 ;
        RECT 178.800 153.000 179.600 153.200 ;
        RECT 183.400 153.000 184.200 153.200 ;
        RECT 178.800 152.400 184.200 153.000 ;
        RECT 184.800 153.000 187.000 153.600 ;
        RECT 184.800 151.800 185.400 153.000 ;
        RECT 186.200 152.800 187.000 153.000 ;
        RECT 188.600 153.200 190.000 154.000 ;
        RECT 188.600 152.200 189.200 153.200 ;
        RECT 180.600 151.400 185.400 151.800 ;
        RECT 175.600 151.200 185.400 151.400 ;
        RECT 186.800 151.600 189.200 152.200 ;
        RECT 175.600 151.000 181.400 151.200 ;
        RECT 175.600 150.800 181.200 151.000 ;
        RECT 158.200 149.800 159.000 150.000 ;
        RECT 158.200 149.200 162.000 149.800 ;
        RECT 162.800 149.600 163.600 150.400 ;
        RECT 166.000 150.300 166.800 150.400 ;
        RECT 167.600 150.300 168.400 150.400 ;
        RECT 166.000 150.200 168.400 150.300 ;
        RECT 182.000 150.200 182.800 150.400 ;
        RECT 166.000 149.700 172.600 150.200 ;
        RECT 166.000 149.600 166.800 149.700 ;
        RECT 167.600 149.600 172.600 149.700 ;
        RECT 161.200 149.000 162.000 149.200 ;
        RECT 163.000 148.400 163.600 149.600 ;
        RECT 171.800 149.400 172.600 149.600 ;
        RECT 177.800 149.600 182.800 150.200 ;
        RECT 177.800 149.400 178.600 149.600 ;
        RECT 180.400 149.400 181.200 149.600 ;
        RECT 170.200 148.400 171.000 148.600 ;
        RECT 179.400 148.400 180.200 148.600 ;
        RECT 186.800 148.400 187.400 151.600 ;
        RECT 193.200 151.200 194.000 159.800 ;
        RECT 189.800 150.600 194.000 151.200 ;
        RECT 189.800 150.400 190.600 150.600 ;
        RECT 191.400 149.800 192.200 150.000 ;
        RECT 188.400 149.200 192.200 149.800 ;
        RECT 188.400 149.000 189.200 149.200 ;
        RECT 163.000 148.300 174.000 148.400 ;
        RECT 176.400 148.300 187.400 148.400 ;
        RECT 163.000 147.800 187.400 148.300 ;
        RECT 163.400 147.600 164.200 147.800 ;
        RECT 156.400 146.600 160.200 147.200 ;
        RECT 154.800 144.800 155.600 146.400 ;
        RECT 153.200 142.200 154.000 144.200 ;
        RECT 156.400 142.200 157.200 146.600 ;
        RECT 159.400 146.400 160.200 146.600 ;
        RECT 169.200 145.600 169.800 147.800 ;
        RECT 172.400 147.700 178.000 147.800 ;
        RECT 172.400 147.600 174.000 147.700 ;
        RECT 176.400 147.600 178.000 147.700 ;
        RECT 167.400 145.400 168.200 145.600 ;
        RECT 161.200 144.200 162.000 145.000 ;
        RECT 165.400 144.800 168.200 145.400 ;
        RECT 169.200 144.800 170.000 145.600 ;
        RECT 165.400 144.200 166.000 144.800 ;
        RECT 170.800 144.200 171.600 145.000 ;
        RECT 160.600 143.600 162.000 144.200 ;
        RECT 160.600 142.200 161.800 143.600 ;
        RECT 165.200 142.200 166.000 144.200 ;
        RECT 169.600 143.600 171.600 144.200 ;
        RECT 169.600 142.200 170.400 143.600 ;
        RECT 174.000 142.200 174.800 147.000 ;
        RECT 175.600 142.200 176.400 147.000 ;
        RECT 180.600 145.600 181.200 147.800 ;
        RECT 186.200 147.600 187.000 147.800 ;
        RECT 193.200 147.200 194.000 150.600 ;
        RECT 190.200 146.600 194.000 147.200 ;
        RECT 190.200 146.400 191.000 146.600 ;
        RECT 178.800 144.200 179.600 145.000 ;
        RECT 180.400 144.800 181.200 145.600 ;
        RECT 182.200 145.400 183.000 145.600 ;
        RECT 182.200 144.800 185.000 145.400 ;
        RECT 184.400 144.200 185.000 144.800 ;
        RECT 188.400 144.200 189.200 145.000 ;
        RECT 178.800 143.600 180.800 144.200 ;
        RECT 180.000 142.200 180.800 143.600 ;
        RECT 184.400 142.200 185.200 144.200 ;
        RECT 188.400 143.600 189.800 144.200 ;
        RECT 188.600 142.200 189.800 143.600 ;
        RECT 193.200 142.200 194.000 146.600 ;
        RECT 4.400 135.200 5.200 139.800 ;
        RECT 9.200 135.200 10.000 139.800 ;
        RECT 3.000 134.600 5.200 135.200 ;
        RECT 7.800 134.600 10.000 135.200 ;
        RECT 14.000 135.800 14.800 139.800 ;
        RECT 15.400 136.400 16.200 137.200 ;
        RECT 3.000 131.600 3.600 134.600 ;
        RECT 4.400 131.600 5.200 133.200 ;
        RECT 7.800 131.600 8.400 134.600 ;
        RECT 9.200 131.600 10.000 133.200 ;
        RECT 12.400 132.800 13.200 134.400 ;
        RECT 10.800 132.200 11.600 132.400 ;
        RECT 14.000 132.200 14.600 135.800 ;
        RECT 15.600 135.600 16.400 136.400 ;
        RECT 17.200 136.000 18.000 139.800 ;
        RECT 20.400 136.000 21.200 139.800 ;
        RECT 17.200 135.800 21.200 136.000 ;
        RECT 22.000 135.800 22.800 139.800 ;
        RECT 17.400 135.400 21.000 135.800 ;
        RECT 18.000 134.400 18.800 134.800 ;
        RECT 22.000 134.400 22.600 135.800 ;
        RECT 23.600 135.600 24.400 137.200 ;
        RECT 15.600 134.300 16.400 134.400 ;
        RECT 17.200 134.300 18.800 134.400 ;
        RECT 15.600 133.800 18.800 134.300 ;
        RECT 15.600 133.700 18.000 133.800 ;
        RECT 15.600 133.600 16.400 133.700 ;
        RECT 17.200 133.600 18.000 133.700 ;
        RECT 20.200 133.600 22.800 134.400 ;
        RECT 15.600 132.200 16.400 132.400 ;
        RECT 10.800 131.600 12.400 132.200 ;
        RECT 14.000 131.600 16.400 132.200 ;
        RECT 18.800 131.600 19.600 133.200 ;
        RECT 2.400 130.800 3.600 131.600 ;
        RECT 7.200 130.800 8.400 131.600 ;
        RECT 11.600 131.200 12.400 131.600 ;
        RECT 3.000 130.200 3.600 130.800 ;
        RECT 7.800 130.200 8.400 130.800 ;
        RECT 15.600 130.200 16.200 131.600 ;
        RECT 20.200 130.200 20.800 133.600 ;
        RECT 22.000 130.200 22.800 130.400 ;
        RECT 3.000 129.600 5.200 130.200 ;
        RECT 7.800 129.600 10.000 130.200 ;
        RECT 4.400 122.200 5.200 129.600 ;
        RECT 9.200 122.200 10.000 129.600 ;
        RECT 10.800 129.600 14.800 130.200 ;
        RECT 10.800 122.200 11.600 129.600 ;
        RECT 14.000 122.200 14.800 129.600 ;
        RECT 15.600 122.200 16.400 130.200 ;
        RECT 19.800 129.600 20.800 130.200 ;
        RECT 21.400 129.600 22.800 130.200 ;
        RECT 19.800 122.200 20.600 129.600 ;
        RECT 21.400 128.400 22.000 129.600 ;
        RECT 21.200 127.600 22.000 128.400 ;
        RECT 25.200 122.200 26.000 139.800 ;
        RECT 29.400 136.400 30.200 139.800 ;
        RECT 28.400 135.800 30.200 136.400 ;
        RECT 31.600 135.800 32.400 139.800 ;
        RECT 34.800 137.800 35.600 139.800 ;
        RECT 26.800 133.600 27.600 135.200 ;
        RECT 28.400 122.200 29.200 135.800 ;
        RECT 31.600 132.400 32.200 135.800 ;
        RECT 34.800 135.600 35.400 137.800 ;
        RECT 36.400 135.600 37.200 137.200 ;
        RECT 41.200 135.800 42.000 139.800 ;
        RECT 46.000 137.800 46.800 139.800 ;
        RECT 33.000 135.000 35.400 135.600 ;
        RECT 31.600 131.600 32.400 132.400 ;
        RECT 33.000 132.000 33.600 135.000 ;
        RECT 34.600 134.300 35.600 134.400 ;
        RECT 39.600 134.300 40.400 134.400 ;
        RECT 34.600 133.700 40.400 134.300 ;
        RECT 34.600 133.600 35.600 133.700 ;
        RECT 34.400 132.800 35.200 133.600 ;
        RECT 39.600 132.800 40.400 133.700 ;
        RECT 38.000 132.200 38.800 132.400 ;
        RECT 41.200 132.200 41.800 135.800 ;
        RECT 46.000 134.400 46.600 137.800 ;
        RECT 47.600 135.600 48.400 137.200 ;
        RECT 46.000 133.600 46.800 134.400 ;
        RECT 42.800 132.200 43.600 132.400 ;
        RECT 30.000 128.800 30.800 130.400 ;
        RECT 31.600 130.200 32.200 131.600 ;
        RECT 33.000 131.400 33.800 132.000 ;
        RECT 38.000 131.600 39.600 132.200 ;
        RECT 41.200 131.600 43.600 132.200 ;
        RECT 33.000 131.200 37.200 131.400 ;
        RECT 38.800 131.200 39.600 131.600 ;
        RECT 33.200 130.800 37.200 131.200 ;
        RECT 31.600 129.600 33.000 130.200 ;
        RECT 32.200 122.200 33.000 129.600 ;
        RECT 36.400 122.200 37.200 130.800 ;
        RECT 42.800 130.200 43.400 131.600 ;
        RECT 44.400 130.800 45.200 132.400 ;
        RECT 46.000 130.200 46.600 133.600 ;
        RECT 38.000 129.600 42.000 130.200 ;
        RECT 38.000 122.200 38.800 129.600 ;
        RECT 41.200 122.200 42.000 129.600 ;
        RECT 42.800 122.200 43.600 130.200 ;
        RECT 45.000 129.400 46.800 130.200 ;
        RECT 45.000 126.400 45.800 129.400 ;
        RECT 45.000 125.600 46.800 126.400 ;
        RECT 45.000 122.200 45.800 125.600 ;
        RECT 49.200 122.200 50.000 139.800 ;
        RECT 50.800 135.600 51.600 137.200 ;
        RECT 60.400 135.800 61.200 139.800 ;
        RECT 64.200 138.400 65.000 139.800 ;
        RECT 64.200 137.600 66.000 138.400 ;
        RECT 61.800 136.400 62.600 137.200 ;
        RECT 64.200 136.400 65.000 137.600 ;
        RECT 58.800 132.800 59.600 134.400 ;
        RECT 57.200 132.200 58.000 132.400 ;
        RECT 60.400 132.200 61.000 135.800 ;
        RECT 62.000 135.600 62.800 136.400 ;
        RECT 64.200 135.800 66.000 136.400 ;
        RECT 68.400 135.800 69.200 139.800 ;
        RECT 70.000 136.000 70.800 139.800 ;
        RECT 73.200 136.000 74.000 139.800 ;
        RECT 70.000 135.800 74.000 136.000 ;
        RECT 76.400 137.800 77.200 139.800 ;
        RECT 62.000 132.300 62.800 132.400 ;
        RECT 63.600 132.300 64.400 132.400 ;
        RECT 62.000 132.200 64.400 132.300 ;
        RECT 57.200 131.600 58.800 132.200 ;
        RECT 60.400 131.700 64.400 132.200 ;
        RECT 60.400 131.600 62.800 131.700 ;
        RECT 63.600 131.600 64.400 131.700 ;
        RECT 58.000 131.200 58.800 131.600 ;
        RECT 62.000 130.200 62.600 131.600 ;
        RECT 57.200 129.600 61.200 130.200 ;
        RECT 57.200 122.200 58.000 129.600 ;
        RECT 60.400 122.200 61.200 129.600 ;
        RECT 62.000 122.200 62.800 130.200 ;
        RECT 63.600 128.800 64.400 130.400 ;
        RECT 65.200 122.200 66.000 135.800 ;
        RECT 66.800 133.600 67.600 135.200 ;
        RECT 68.600 134.400 69.200 135.800 ;
        RECT 70.200 135.400 73.800 135.800 ;
        RECT 72.400 134.400 73.200 134.800 ;
        RECT 76.400 134.400 77.000 137.800 ;
        RECT 78.000 136.300 78.800 137.200 ;
        RECT 80.200 136.400 81.000 139.800 ;
        RECT 80.200 136.300 82.000 136.400 ;
        RECT 78.000 135.700 82.000 136.300 ;
        RECT 78.000 135.600 78.800 135.700 ;
        RECT 68.400 133.600 71.000 134.400 ;
        RECT 72.400 134.300 74.000 134.400 ;
        RECT 74.800 134.300 75.600 134.400 ;
        RECT 72.400 133.800 75.600 134.300 ;
        RECT 73.200 133.700 75.600 133.800 ;
        RECT 73.200 133.600 74.000 133.700 ;
        RECT 74.800 133.600 75.600 133.700 ;
        RECT 76.400 133.600 77.200 134.400 ;
        RECT 68.400 130.200 69.200 130.400 ;
        RECT 70.400 130.200 71.000 133.600 ;
        RECT 71.600 131.600 72.400 133.200 ;
        RECT 73.200 132.300 74.000 132.400 ;
        RECT 74.800 132.300 75.600 132.400 ;
        RECT 73.200 131.700 75.600 132.300 ;
        RECT 73.200 131.600 74.000 131.700 ;
        RECT 74.800 130.800 75.600 131.700 ;
        RECT 76.400 132.300 77.000 133.600 ;
        RECT 79.600 132.300 80.400 132.400 ;
        RECT 76.400 131.700 80.400 132.300 ;
        RECT 76.400 130.200 77.000 131.700 ;
        RECT 79.600 131.600 80.400 131.700 ;
        RECT 68.400 129.600 69.800 130.200 ;
        RECT 70.400 129.600 71.400 130.200 ;
        RECT 69.200 128.400 69.800 129.600 ;
        RECT 69.200 127.600 70.000 128.400 ;
        RECT 70.600 122.200 71.400 129.600 ;
        RECT 75.400 129.400 77.200 130.200 ;
        RECT 75.400 122.200 76.200 129.400 ;
        RECT 79.600 128.800 80.400 130.400 ;
        RECT 81.200 122.200 82.000 135.700 ;
        RECT 84.400 135.400 85.200 139.800 ;
        RECT 88.600 138.400 89.800 139.800 ;
        RECT 88.600 137.800 90.000 138.400 ;
        RECT 93.200 137.800 94.000 139.800 ;
        RECT 97.600 138.400 98.400 139.800 ;
        RECT 97.600 137.800 99.600 138.400 ;
        RECT 89.200 137.000 90.000 137.800 ;
        RECT 93.400 137.200 94.000 137.800 ;
        RECT 93.400 136.600 96.200 137.200 ;
        RECT 95.400 136.400 96.200 136.600 ;
        RECT 97.200 136.400 98.000 137.200 ;
        RECT 98.800 137.000 99.600 137.800 ;
        RECT 87.400 135.400 88.200 135.600 ;
        RECT 82.800 133.600 83.600 135.200 ;
        RECT 84.400 134.800 88.200 135.400 ;
        RECT 84.400 131.400 85.200 134.800 ;
        RECT 91.400 134.200 92.200 134.400 ;
        RECT 97.200 134.200 97.800 136.400 ;
        RECT 102.000 135.000 102.800 139.800 ;
        RECT 103.600 135.400 104.400 139.800 ;
        RECT 107.800 138.400 109.000 139.800 ;
        RECT 107.800 137.800 109.200 138.400 ;
        RECT 112.400 137.800 113.200 139.800 ;
        RECT 116.800 138.400 117.600 139.800 ;
        RECT 116.800 137.800 118.800 138.400 ;
        RECT 108.400 137.000 109.200 137.800 ;
        RECT 112.600 137.200 113.200 137.800 ;
        RECT 112.600 136.600 115.400 137.200 ;
        RECT 114.600 136.400 115.400 136.600 ;
        RECT 116.400 136.400 117.200 137.200 ;
        RECT 118.000 137.000 118.800 137.800 ;
        RECT 106.600 135.400 107.400 135.600 ;
        RECT 103.600 134.800 107.400 135.400 ;
        RECT 100.400 134.200 102.000 134.400 ;
        RECT 91.000 133.600 102.000 134.200 ;
        RECT 89.200 132.800 90.000 133.000 ;
        RECT 86.200 132.200 90.000 132.800 ;
        RECT 86.200 132.000 87.000 132.200 ;
        RECT 87.800 131.400 88.600 131.600 ;
        RECT 84.400 130.800 88.600 131.400 ;
        RECT 84.400 122.200 85.200 130.800 ;
        RECT 91.000 130.400 91.600 133.600 ;
        RECT 98.200 133.400 99.000 133.600 ;
        RECT 99.800 132.400 100.600 132.600 ;
        RECT 95.600 131.800 100.600 132.400 ;
        RECT 95.600 131.600 96.400 131.800 ;
        RECT 103.600 131.400 104.400 134.800 ;
        RECT 105.200 133.600 106.000 134.800 ;
        RECT 110.600 134.200 111.400 134.400 ;
        RECT 116.400 134.200 117.000 136.400 ;
        RECT 121.200 135.000 122.000 139.800 ;
        RECT 124.400 137.800 125.200 139.800 ;
        RECT 122.800 135.600 123.600 137.200 ;
        RECT 124.600 134.400 125.200 137.800 ;
        RECT 128.200 136.400 129.000 139.800 ;
        RECT 132.600 136.400 133.400 137.200 ;
        RECT 128.200 135.800 130.000 136.400 ;
        RECT 119.600 134.200 121.200 134.400 ;
        RECT 110.200 133.600 121.200 134.200 ;
        RECT 124.400 133.600 125.200 134.400 ;
        RECT 108.400 132.800 109.200 133.000 ;
        RECT 105.400 132.200 109.200 132.800 ;
        RECT 110.200 132.400 110.800 133.600 ;
        RECT 117.400 133.400 118.200 133.600 ;
        RECT 119.000 132.400 119.800 132.600 ;
        RECT 105.400 132.000 106.200 132.200 ;
        RECT 110.000 131.600 110.800 132.400 ;
        RECT 114.800 131.800 119.800 132.400 ;
        RECT 122.800 132.300 123.600 132.400 ;
        RECT 124.600 132.300 125.200 133.600 ;
        RECT 114.800 131.600 115.600 131.800 ;
        RECT 122.800 131.700 125.200 132.300 ;
        RECT 122.800 131.600 123.600 131.700 ;
        RECT 107.000 131.400 107.800 131.600 ;
        RECT 97.200 131.000 102.800 131.200 ;
        RECT 97.000 130.800 102.800 131.000 ;
        RECT 89.200 129.800 91.600 130.400 ;
        RECT 93.000 130.600 102.800 130.800 ;
        RECT 93.000 130.200 97.800 130.600 ;
        RECT 89.200 128.800 89.800 129.800 ;
        RECT 88.400 128.000 89.800 128.800 ;
        RECT 91.400 129.000 92.200 129.200 ;
        RECT 93.000 129.000 93.600 130.200 ;
        RECT 91.400 128.400 93.600 129.000 ;
        RECT 94.200 129.000 99.600 129.600 ;
        RECT 94.200 128.800 95.000 129.000 ;
        RECT 98.800 128.800 99.600 129.000 ;
        RECT 92.600 127.400 93.400 127.600 ;
        RECT 95.400 127.400 96.200 127.600 ;
        RECT 89.200 126.200 90.000 127.000 ;
        RECT 92.600 126.800 96.200 127.400 ;
        RECT 93.400 126.200 94.000 126.800 ;
        RECT 98.800 126.200 99.600 127.000 ;
        RECT 88.600 122.200 89.800 126.200 ;
        RECT 93.200 122.200 94.000 126.200 ;
        RECT 97.600 125.600 99.600 126.200 ;
        RECT 97.600 122.200 98.400 125.600 ;
        RECT 102.000 122.200 102.800 130.600 ;
        RECT 103.600 130.800 107.800 131.400 ;
        RECT 103.600 122.200 104.400 130.800 ;
        RECT 110.200 130.400 110.800 131.600 ;
        RECT 116.400 131.000 122.000 131.200 ;
        RECT 116.200 130.800 122.000 131.000 ;
        RECT 108.400 129.800 110.800 130.400 ;
        RECT 112.200 130.600 122.000 130.800 ;
        RECT 112.200 130.200 117.000 130.600 ;
        RECT 108.400 128.800 109.000 129.800 ;
        RECT 107.600 128.000 109.000 128.800 ;
        RECT 110.600 129.000 111.400 129.200 ;
        RECT 112.200 129.000 112.800 130.200 ;
        RECT 110.600 128.400 112.800 129.000 ;
        RECT 113.400 129.000 118.800 129.600 ;
        RECT 113.400 128.800 114.200 129.000 ;
        RECT 118.000 128.800 118.800 129.000 ;
        RECT 111.800 127.400 112.600 127.600 ;
        RECT 114.600 127.400 115.400 127.600 ;
        RECT 108.400 126.200 109.200 127.000 ;
        RECT 111.800 126.800 115.400 127.400 ;
        RECT 112.600 126.200 113.200 126.800 ;
        RECT 118.000 126.200 118.800 127.000 ;
        RECT 107.800 122.200 109.000 126.200 ;
        RECT 112.400 122.200 113.200 126.200 ;
        RECT 116.800 125.600 118.800 126.200 ;
        RECT 116.800 122.200 117.600 125.600 ;
        RECT 121.200 122.200 122.000 130.600 ;
        RECT 124.600 130.200 125.200 131.700 ;
        RECT 126.000 130.800 126.800 132.400 ;
        RECT 124.400 129.400 126.200 130.200 ;
        RECT 125.400 122.200 126.200 129.400 ;
        RECT 127.600 128.800 128.400 130.400 ;
        RECT 129.200 122.200 130.000 135.800 ;
        RECT 132.400 135.600 133.200 136.400 ;
        RECT 134.000 135.800 134.800 139.800 ;
        RECT 130.800 133.600 131.600 135.200 ;
        RECT 132.400 132.200 133.200 132.400 ;
        RECT 134.200 132.200 134.800 135.800 ;
        RECT 143.600 135.600 144.400 137.200 ;
        RECT 135.600 132.800 136.400 134.400 ;
        RECT 137.200 132.200 138.000 132.400 ;
        RECT 132.400 131.600 134.800 132.200 ;
        RECT 136.400 131.600 138.000 132.200 ;
        RECT 132.600 130.200 133.200 131.600 ;
        RECT 136.400 131.200 137.200 131.600 ;
        RECT 130.800 128.300 131.600 128.400 ;
        RECT 132.400 128.300 133.200 130.200 ;
        RECT 130.800 127.700 133.200 128.300 ;
        RECT 130.800 127.600 131.600 127.700 ;
        RECT 132.400 122.200 133.200 127.700 ;
        RECT 134.000 129.600 138.000 130.200 ;
        RECT 134.000 122.200 134.800 129.600 ;
        RECT 137.200 122.200 138.000 129.600 ;
        RECT 145.200 122.200 146.000 139.800 ;
        RECT 148.400 137.800 149.200 139.800 ;
        RECT 146.800 135.600 147.600 137.200 ;
        RECT 148.600 134.400 149.200 137.800 ;
        RECT 154.800 135.800 155.600 139.800 ;
        RECT 156.200 136.400 157.000 137.200 ;
        RECT 148.400 134.300 149.200 134.400 ;
        RECT 153.200 134.300 154.000 134.400 ;
        RECT 148.400 133.700 154.000 134.300 ;
        RECT 148.400 133.600 149.200 133.700 ;
        RECT 148.600 130.200 149.200 133.600 ;
        RECT 153.200 132.800 154.000 133.700 ;
        RECT 150.000 130.800 150.800 132.400 ;
        RECT 151.600 132.200 152.400 132.400 ;
        RECT 154.800 132.200 155.400 135.800 ;
        RECT 156.400 135.600 157.200 136.400 ;
        RECT 158.000 136.000 158.800 139.800 ;
        RECT 161.200 136.000 162.000 139.800 ;
        RECT 158.000 135.800 162.000 136.000 ;
        RECT 162.800 135.800 163.600 139.800 ;
        RECT 167.000 136.400 167.800 139.800 ;
        RECT 169.400 136.400 170.200 137.200 ;
        RECT 166.000 136.300 167.800 136.400 ;
        RECT 169.200 136.300 170.000 136.400 ;
        RECT 158.200 135.400 161.800 135.800 ;
        RECT 158.800 134.400 159.600 134.800 ;
        RECT 162.800 134.400 163.400 135.800 ;
        RECT 166.000 135.700 170.000 136.300 ;
        RECT 170.800 135.800 171.600 139.800 ;
        RECT 156.400 134.300 157.200 134.400 ;
        RECT 158.000 134.300 159.600 134.400 ;
        RECT 156.400 133.800 159.600 134.300 ;
        RECT 156.400 133.700 158.800 133.800 ;
        RECT 156.400 133.600 157.200 133.700 ;
        RECT 158.000 133.600 158.800 133.700 ;
        RECT 161.000 133.600 163.600 134.400 ;
        RECT 164.400 133.600 165.200 135.200 ;
        RECT 156.400 132.200 157.200 132.400 ;
        RECT 151.600 131.600 153.200 132.200 ;
        RECT 154.800 131.600 157.200 132.200 ;
        RECT 159.600 131.600 160.400 133.200 ;
        RECT 152.400 131.200 153.200 131.600 ;
        RECT 156.400 130.200 157.000 131.600 ;
        RECT 161.000 130.200 161.600 133.600 ;
        RECT 162.800 130.200 163.600 130.400 ;
        RECT 148.400 129.400 150.200 130.200 ;
        RECT 149.400 122.200 150.200 129.400 ;
        RECT 151.600 129.600 155.600 130.200 ;
        RECT 151.600 122.200 152.400 129.600 ;
        RECT 154.800 122.200 155.600 129.600 ;
        RECT 156.400 122.200 157.200 130.200 ;
        RECT 160.600 129.600 161.600 130.200 ;
        RECT 162.200 129.600 163.600 130.200 ;
        RECT 160.600 122.200 161.400 129.600 ;
        RECT 162.200 128.400 162.800 129.600 ;
        RECT 162.000 127.600 162.800 128.400 ;
        RECT 166.000 122.200 166.800 135.700 ;
        RECT 169.200 135.600 170.000 135.700 ;
        RECT 169.200 132.200 170.000 132.400 ;
        RECT 171.000 132.200 171.600 135.800 ;
        RECT 175.600 135.000 176.400 139.800 ;
        RECT 180.000 138.400 180.800 139.800 ;
        RECT 178.800 137.800 180.800 138.400 ;
        RECT 184.400 137.800 185.200 139.800 ;
        RECT 188.600 138.400 189.800 139.800 ;
        RECT 188.400 137.800 189.800 138.400 ;
        RECT 178.800 137.000 179.600 137.800 ;
        RECT 184.400 137.200 185.000 137.800 ;
        RECT 180.400 136.400 181.200 137.200 ;
        RECT 182.200 136.600 185.000 137.200 ;
        RECT 188.400 137.000 189.200 137.800 ;
        RECT 182.200 136.400 183.000 136.600 ;
        RECT 172.400 132.800 173.200 134.400 ;
        RECT 176.400 134.200 178.000 134.400 ;
        RECT 180.600 134.200 181.200 136.400 ;
        RECT 190.200 135.400 191.000 135.600 ;
        RECT 193.200 135.400 194.000 139.800 ;
        RECT 190.200 134.800 194.000 135.400 ;
        RECT 186.200 134.200 187.000 134.400 ;
        RECT 176.400 133.600 187.400 134.200 ;
        RECT 179.400 133.400 180.200 133.600 ;
        RECT 177.800 132.400 178.600 132.600 ;
        RECT 174.000 132.200 174.800 132.400 ;
        RECT 169.200 131.600 171.600 132.200 ;
        RECT 173.200 131.600 174.800 132.200 ;
        RECT 177.800 132.300 182.800 132.400 ;
        RECT 183.600 132.300 184.400 132.400 ;
        RECT 177.800 131.800 184.400 132.300 ;
        RECT 182.000 131.700 184.400 131.800 ;
        RECT 182.000 131.600 182.800 131.700 ;
        RECT 183.600 131.600 184.400 131.700 ;
        RECT 167.600 128.800 168.400 130.400 ;
        RECT 169.400 130.200 170.000 131.600 ;
        RECT 173.200 131.200 174.000 131.600 ;
        RECT 175.600 131.000 181.200 131.200 ;
        RECT 175.600 130.800 181.400 131.000 ;
        RECT 175.600 130.600 185.400 130.800 ;
        RECT 169.200 122.200 170.000 130.200 ;
        RECT 170.800 129.600 174.800 130.200 ;
        RECT 170.800 122.200 171.600 129.600 ;
        RECT 174.000 122.200 174.800 129.600 ;
        RECT 175.600 122.200 176.400 130.600 ;
        RECT 180.600 130.200 185.400 130.600 ;
        RECT 178.800 129.000 184.200 129.600 ;
        RECT 178.800 128.800 179.600 129.000 ;
        RECT 183.400 128.800 184.200 129.000 ;
        RECT 184.800 129.000 185.400 130.200 ;
        RECT 186.800 130.400 187.400 133.600 ;
        RECT 188.400 132.800 189.200 133.000 ;
        RECT 188.400 132.200 192.200 132.800 ;
        RECT 191.400 132.000 192.200 132.200 ;
        RECT 189.800 131.400 190.600 131.600 ;
        RECT 193.200 131.400 194.000 134.800 ;
        RECT 189.800 130.800 194.000 131.400 ;
        RECT 186.800 129.800 189.200 130.400 ;
        RECT 186.200 129.000 187.000 129.200 ;
        RECT 184.800 128.400 187.000 129.000 ;
        RECT 188.600 128.800 189.200 129.800 ;
        RECT 188.600 128.000 190.000 128.800 ;
        RECT 182.200 127.400 183.000 127.600 ;
        RECT 185.000 127.400 185.800 127.600 ;
        RECT 178.800 126.200 179.600 127.000 ;
        RECT 182.200 126.800 185.800 127.400 ;
        RECT 184.400 126.200 185.000 126.800 ;
        RECT 188.400 126.200 189.200 127.000 ;
        RECT 178.800 125.600 180.800 126.200 ;
        RECT 180.000 122.200 180.800 125.600 ;
        RECT 184.400 122.200 185.200 126.200 ;
        RECT 188.600 122.200 189.800 126.200 ;
        RECT 193.200 122.200 194.000 130.800 ;
        RECT 4.400 112.400 5.200 119.800 ;
        RECT 3.000 111.800 5.200 112.400 ;
        RECT 3.000 111.200 3.600 111.800 ;
        RECT 2.400 110.400 3.600 111.200 ;
        RECT 6.000 111.200 6.800 119.800 ;
        RECT 10.200 115.800 11.400 119.800 ;
        RECT 14.800 115.800 15.600 119.800 ;
        RECT 19.200 116.400 20.000 119.800 ;
        RECT 19.200 115.800 21.200 116.400 ;
        RECT 10.800 115.000 11.600 115.800 ;
        RECT 15.000 115.200 15.600 115.800 ;
        RECT 14.200 114.600 17.800 115.200 ;
        RECT 20.400 115.000 21.200 115.800 ;
        RECT 14.200 114.400 15.000 114.600 ;
        RECT 17.000 114.400 17.800 114.600 ;
        RECT 10.000 113.200 11.400 114.000 ;
        RECT 10.800 112.200 11.400 113.200 ;
        RECT 13.000 113.000 15.200 113.600 ;
        RECT 13.000 112.800 13.800 113.000 ;
        RECT 10.800 111.600 13.200 112.200 ;
        RECT 6.000 110.600 10.200 111.200 ;
        RECT 3.000 107.400 3.600 110.400 ;
        RECT 4.400 108.800 5.200 110.400 ;
        RECT 3.000 106.800 5.200 107.400 ;
        RECT 4.400 102.200 5.200 106.800 ;
        RECT 6.000 107.200 6.800 110.600 ;
        RECT 9.400 110.400 10.200 110.600 ;
        RECT 7.800 109.800 8.600 110.000 ;
        RECT 7.800 109.200 11.600 109.800 ;
        RECT 10.800 109.000 11.600 109.200 ;
        RECT 12.600 108.400 13.200 111.600 ;
        RECT 14.600 111.800 15.200 113.000 ;
        RECT 15.800 113.000 16.600 113.200 ;
        RECT 20.400 113.000 21.200 113.200 ;
        RECT 15.800 112.400 21.200 113.000 ;
        RECT 14.600 111.400 19.400 111.800 ;
        RECT 23.600 111.400 24.400 119.800 ;
        RECT 14.600 111.200 24.400 111.400 ;
        RECT 18.600 111.000 24.400 111.200 ;
        RECT 18.800 110.800 24.400 111.000 ;
        RECT 25.200 111.600 26.000 119.800 ;
        RECT 28.400 115.800 29.200 119.800 ;
        RECT 28.400 111.600 29.000 115.800 ;
        RECT 25.200 110.400 25.800 111.600 ;
        RECT 26.600 111.000 29.000 111.600 ;
        RECT 17.200 110.200 18.000 110.400 ;
        RECT 17.200 109.600 22.200 110.200 ;
        RECT 18.800 109.400 19.600 109.600 ;
        RECT 21.400 109.400 22.200 109.600 ;
        RECT 25.200 109.600 26.000 110.400 ;
        RECT 19.800 108.400 20.600 108.600 ;
        RECT 12.600 107.800 23.600 108.400 ;
        RECT 13.000 107.600 13.800 107.800 ;
        RECT 17.200 107.600 18.000 107.800 ;
        RECT 6.000 106.600 9.800 107.200 ;
        RECT 6.000 102.200 6.800 106.600 ;
        RECT 9.000 106.400 9.800 106.600 ;
        RECT 18.800 105.600 19.400 107.800 ;
        RECT 22.000 107.600 23.600 107.800 ;
        RECT 17.000 105.400 17.800 105.600 ;
        RECT 10.800 104.200 11.600 105.000 ;
        RECT 15.000 104.800 17.800 105.400 ;
        RECT 18.800 104.800 19.600 105.600 ;
        RECT 15.000 104.200 15.600 104.800 ;
        RECT 20.400 104.200 21.200 105.000 ;
        RECT 10.200 103.600 11.600 104.200 ;
        RECT 10.200 102.200 11.400 103.600 ;
        RECT 14.800 102.200 15.600 104.200 ;
        RECT 19.200 103.600 21.200 104.200 ;
        RECT 19.200 102.200 20.000 103.600 ;
        RECT 23.600 102.200 24.400 107.000 ;
        RECT 25.200 106.200 25.800 109.600 ;
        RECT 26.600 107.600 27.200 111.000 ;
        RECT 28.400 109.600 29.200 110.400 ;
        RECT 28.400 108.800 29.000 109.600 ;
        RECT 28.000 108.200 29.000 108.800 ;
        RECT 28.000 108.000 28.800 108.200 ;
        RECT 30.000 107.600 30.800 109.200 ;
        RECT 26.400 107.400 27.200 107.600 ;
        RECT 26.400 107.000 29.400 107.400 ;
        RECT 26.400 106.800 30.600 107.000 ;
        RECT 28.800 106.400 30.600 106.800 ;
        RECT 30.000 106.200 30.600 106.400 ;
        RECT 33.200 106.300 34.000 119.800 ;
        RECT 37.400 118.400 38.200 119.800 ;
        RECT 42.200 118.400 43.000 119.800 ;
        RECT 36.400 117.600 38.200 118.400 ;
        RECT 41.200 117.600 43.000 118.400 ;
        RECT 37.400 112.600 38.200 117.600 ;
        RECT 36.400 111.800 38.200 112.600 ;
        RECT 42.200 112.400 43.000 117.600 ;
        RECT 46.000 115.800 46.800 119.800 ;
        RECT 46.200 115.600 46.800 115.800 ;
        RECT 49.200 115.800 50.000 119.800 ;
        RECT 57.200 115.800 58.000 119.800 ;
        RECT 49.200 115.600 49.800 115.800 ;
        RECT 46.200 115.000 49.800 115.600 ;
        RECT 57.400 115.600 58.000 115.800 ;
        RECT 60.400 115.800 61.200 119.800 ;
        RECT 65.200 115.800 66.000 119.800 ;
        RECT 60.400 115.600 61.000 115.800 ;
        RECT 57.400 115.000 61.000 115.600 ;
        RECT 43.600 113.600 44.400 114.400 ;
        RECT 43.800 112.400 44.400 113.600 ;
        RECT 46.200 112.400 46.800 115.000 ;
        RECT 47.600 112.800 48.400 114.400 ;
        RECT 57.400 112.400 58.000 115.000 ;
        RECT 58.800 112.800 59.600 114.400 ;
        RECT 42.200 111.800 43.200 112.400 ;
        RECT 43.800 111.800 45.200 112.400 ;
        RECT 36.600 108.400 37.200 111.800 ;
        RECT 38.000 110.300 38.800 111.200 ;
        RECT 41.200 110.300 42.000 110.400 ;
        RECT 38.000 109.700 42.000 110.300 ;
        RECT 38.000 109.600 38.800 109.700 ;
        RECT 41.200 108.800 42.000 109.700 ;
        RECT 42.600 108.400 43.200 111.800 ;
        RECT 44.400 111.600 45.200 111.800 ;
        RECT 46.000 111.600 46.800 112.400 ;
        RECT 46.200 108.400 46.800 111.600 ;
        RECT 50.800 110.800 51.600 112.400 ;
        RECT 57.200 111.600 58.000 112.400 ;
        RECT 48.400 109.600 50.000 110.400 ;
        RECT 57.400 108.400 58.000 111.600 ;
        RECT 62.000 112.300 62.800 112.400 ;
        RECT 63.600 112.300 64.400 112.400 ;
        RECT 62.000 111.700 64.400 112.300 ;
        RECT 62.000 110.800 62.800 111.700 ;
        RECT 63.600 111.600 64.400 111.700 ;
        RECT 65.400 111.600 66.000 115.800 ;
        RECT 68.400 112.300 69.200 119.800 ;
        RECT 70.000 112.300 70.800 112.400 ;
        RECT 68.400 111.800 70.800 112.300 ;
        RECT 68.500 111.700 70.800 111.800 ;
        RECT 65.400 111.000 67.800 111.600 ;
        RECT 59.600 109.600 61.200 110.400 ;
        RECT 65.200 109.600 66.000 110.400 ;
        RECT 36.400 107.600 37.200 108.400 ;
        RECT 39.600 108.200 40.400 108.400 ;
        RECT 39.600 107.600 41.200 108.200 ;
        RECT 42.600 107.600 45.200 108.400 ;
        RECT 46.200 108.200 47.800 108.400 ;
        RECT 57.400 108.200 59.000 108.400 ;
        RECT 46.200 107.800 48.000 108.200 ;
        RECT 57.400 107.800 59.200 108.200 ;
        RECT 34.800 106.300 35.600 106.400 ;
        RECT 25.200 105.200 26.600 106.200 ;
        RECT 25.800 102.200 26.600 105.200 ;
        RECT 30.000 102.200 30.800 106.200 ;
        RECT 33.200 105.700 35.600 106.300 ;
        RECT 33.200 102.200 34.000 105.700 ;
        RECT 34.800 104.800 35.600 105.700 ;
        RECT 36.600 104.200 37.200 107.600 ;
        RECT 40.400 107.200 41.200 107.600 ;
        RECT 39.800 106.200 43.400 106.600 ;
        RECT 44.400 106.200 45.000 107.600 ;
        RECT 36.400 102.200 37.200 104.200 ;
        RECT 39.600 106.000 43.600 106.200 ;
        RECT 39.600 102.200 40.400 106.000 ;
        RECT 42.800 102.200 43.600 106.000 ;
        RECT 44.400 102.200 45.200 106.200 ;
        RECT 47.200 102.200 48.000 107.800 ;
        RECT 58.400 102.200 59.200 107.800 ;
        RECT 63.600 107.600 64.400 109.200 ;
        RECT 65.400 108.800 66.000 109.600 ;
        RECT 65.400 108.200 66.400 108.800 ;
        RECT 65.600 108.000 66.400 108.200 ;
        RECT 67.200 107.600 67.800 111.000 ;
        RECT 68.600 110.400 69.200 111.700 ;
        RECT 70.000 111.600 70.800 111.700 ;
        RECT 68.400 109.600 69.200 110.400 ;
        RECT 67.200 107.400 68.000 107.600 ;
        RECT 65.000 107.000 68.000 107.400 ;
        RECT 63.800 106.800 68.000 107.000 ;
        RECT 63.800 106.400 65.600 106.800 ;
        RECT 63.800 106.200 64.400 106.400 ;
        RECT 68.600 106.200 69.200 109.600 ;
        RECT 71.600 110.300 72.400 119.800 ;
        RECT 73.200 111.600 74.000 113.200 ;
        RECT 77.400 112.600 78.200 119.800 ;
        RECT 76.400 111.800 78.200 112.600 ;
        RECT 73.200 110.300 74.000 110.400 ;
        RECT 71.600 109.700 74.000 110.300 ;
        RECT 70.000 106.800 70.800 108.400 ;
        RECT 63.600 102.200 64.400 106.200 ;
        RECT 67.800 105.200 69.200 106.200 ;
        RECT 71.600 106.200 72.400 109.700 ;
        RECT 73.200 109.600 74.000 109.700 ;
        RECT 76.600 108.400 77.200 111.800 ;
        RECT 78.000 109.600 78.800 111.200 ;
        RECT 76.400 107.600 77.200 108.400 ;
        RECT 71.600 105.600 73.400 106.200 ;
        RECT 67.800 102.200 68.600 105.200 ;
        RECT 72.600 102.200 73.400 105.600 ;
        RECT 74.800 104.800 75.600 106.400 ;
        RECT 76.600 104.400 77.200 107.600 ;
        RECT 79.600 106.800 80.400 108.400 ;
        RECT 81.200 106.200 82.000 119.800 ;
        RECT 85.200 113.600 86.000 114.400 ;
        RECT 82.800 111.600 83.600 113.200 ;
        RECT 85.200 112.400 85.800 113.600 ;
        RECT 86.600 112.400 87.400 119.800 ;
        RECT 84.400 111.800 85.800 112.400 ;
        RECT 86.400 111.800 87.400 112.400 ;
        RECT 90.800 111.800 91.600 119.800 ;
        RECT 92.400 112.400 93.200 119.800 ;
        RECT 95.600 112.400 96.400 119.800 ;
        RECT 92.400 111.800 96.400 112.400 ;
        RECT 84.400 111.600 85.200 111.800 ;
        RECT 86.400 108.400 87.000 111.800 ;
        RECT 91.000 110.400 91.600 111.800 ;
        RECT 94.800 110.400 95.600 110.800 ;
        RECT 87.600 108.800 88.400 110.400 ;
        RECT 90.800 109.800 93.200 110.400 ;
        RECT 94.800 110.300 96.400 110.400 ;
        RECT 97.200 110.300 98.000 119.800 ;
        RECT 98.800 114.300 99.600 114.400 ;
        RECT 100.400 114.300 101.200 119.800 ;
        RECT 104.600 115.800 105.800 119.800 ;
        RECT 109.200 115.800 110.000 119.800 ;
        RECT 113.600 116.400 114.400 119.800 ;
        RECT 113.600 115.800 115.600 116.400 ;
        RECT 105.200 115.000 106.000 115.800 ;
        RECT 109.400 115.200 110.000 115.800 ;
        RECT 108.600 114.600 112.200 115.200 ;
        RECT 114.800 115.000 115.600 115.800 ;
        RECT 108.600 114.400 109.400 114.600 ;
        RECT 111.400 114.400 112.200 114.600 ;
        RECT 98.800 113.700 101.200 114.300 ;
        RECT 98.800 113.600 99.600 113.700 ;
        RECT 94.800 109.800 98.000 110.300 ;
        RECT 90.800 109.600 91.600 109.800 ;
        RECT 92.400 109.600 93.200 109.800 ;
        RECT 95.600 109.700 98.000 109.800 ;
        RECT 95.600 109.600 96.400 109.700 ;
        RECT 84.400 107.600 87.000 108.400 ;
        RECT 89.200 108.200 90.000 108.400 ;
        RECT 88.400 107.600 90.000 108.200 ;
        RECT 84.600 106.200 85.200 107.600 ;
        RECT 88.400 107.200 89.200 107.600 ;
        RECT 86.200 106.200 89.800 106.600 ;
        RECT 81.200 105.600 83.000 106.200 ;
        RECT 76.400 102.200 77.200 104.400 ;
        RECT 82.200 104.400 83.000 105.600 ;
        RECT 82.200 103.600 83.600 104.400 ;
        RECT 82.200 102.200 83.000 103.600 ;
        RECT 84.400 102.200 85.200 106.200 ;
        RECT 86.000 106.000 90.000 106.200 ;
        RECT 86.000 102.200 86.800 106.000 ;
        RECT 89.200 102.200 90.000 106.000 ;
        RECT 90.800 105.600 91.600 106.400 ;
        RECT 92.600 106.200 93.200 109.600 ;
        RECT 94.000 107.600 94.800 109.200 ;
        RECT 95.600 108.300 96.400 108.400 ;
        RECT 97.200 108.300 98.000 109.700 ;
        RECT 95.600 107.700 98.000 108.300 ;
        RECT 95.600 107.600 96.400 107.700 ;
        RECT 91.000 104.800 91.800 105.600 ;
        RECT 92.400 102.200 93.200 106.200 ;
        RECT 97.200 102.200 98.000 107.700 ;
        RECT 100.400 111.200 101.200 113.700 ;
        RECT 104.400 113.200 105.800 114.000 ;
        RECT 105.200 112.200 105.800 113.200 ;
        RECT 107.400 113.000 109.600 113.600 ;
        RECT 107.400 112.800 108.200 113.000 ;
        RECT 105.200 111.600 107.600 112.200 ;
        RECT 100.400 110.600 104.600 111.200 ;
        RECT 100.400 107.200 101.200 110.600 ;
        RECT 103.800 110.400 104.600 110.600 ;
        RECT 102.200 109.800 103.000 110.000 ;
        RECT 102.200 109.200 106.000 109.800 ;
        RECT 105.200 109.000 106.000 109.200 ;
        RECT 107.000 108.400 107.600 111.600 ;
        RECT 109.000 111.800 109.600 113.000 ;
        RECT 110.200 113.000 111.000 113.200 ;
        RECT 114.800 113.000 115.600 113.200 ;
        RECT 110.200 112.400 115.600 113.000 ;
        RECT 109.000 111.400 113.800 111.800 ;
        RECT 118.000 111.400 118.800 119.800 ;
        RECT 120.200 112.600 121.000 119.800 ;
        RECT 120.200 111.800 122.000 112.600 ;
        RECT 109.000 111.200 118.800 111.400 ;
        RECT 113.000 111.000 118.800 111.200 ;
        RECT 113.200 110.800 118.800 111.000 ;
        RECT 111.600 110.200 112.400 110.400 ;
        RECT 111.600 109.600 116.600 110.200 ;
        RECT 119.600 109.600 120.400 111.200 ;
        RECT 115.800 109.400 116.600 109.600 ;
        RECT 114.200 108.400 115.000 108.600 ;
        RECT 121.200 108.400 121.800 111.800 ;
        RECT 124.400 111.400 125.200 119.800 ;
        RECT 128.800 116.400 129.600 119.800 ;
        RECT 127.600 115.800 129.600 116.400 ;
        RECT 133.200 115.800 134.000 119.800 ;
        RECT 137.400 115.800 138.600 119.800 ;
        RECT 127.600 115.000 128.400 115.800 ;
        RECT 133.200 115.200 133.800 115.800 ;
        RECT 131.000 114.600 134.600 115.200 ;
        RECT 137.200 115.000 138.000 115.800 ;
        RECT 131.000 114.400 131.800 114.600 ;
        RECT 133.800 114.400 134.600 114.600 ;
        RECT 138.200 114.000 139.600 114.400 ;
        RECT 137.400 113.600 139.600 114.000 ;
        RECT 127.600 113.000 128.400 113.200 ;
        RECT 132.200 113.000 133.000 113.200 ;
        RECT 127.600 112.400 133.000 113.000 ;
        RECT 133.600 113.000 135.800 113.600 ;
        RECT 133.600 111.800 134.200 113.000 ;
        RECT 135.000 112.800 135.800 113.000 ;
        RECT 137.400 113.200 138.800 113.600 ;
        RECT 137.400 112.200 138.000 113.200 ;
        RECT 129.400 111.400 134.200 111.800 ;
        RECT 124.400 111.200 134.200 111.400 ;
        RECT 135.600 111.600 138.000 112.200 ;
        RECT 124.400 111.000 130.200 111.200 ;
        RECT 124.400 110.800 130.000 111.000 ;
        RECT 130.800 110.200 131.600 110.400 ;
        RECT 126.600 109.600 131.600 110.200 ;
        RECT 126.600 109.400 127.400 109.600 ;
        RECT 129.200 109.400 130.000 109.600 ;
        RECT 128.200 108.400 129.000 108.600 ;
        RECT 135.600 108.400 136.200 111.600 ;
        RECT 142.000 111.200 142.800 119.800 ;
        RECT 149.200 113.600 150.000 114.400 ;
        RECT 149.200 112.400 149.800 113.600 ;
        RECT 150.600 112.400 151.400 119.800 ;
        RECT 146.800 112.300 147.600 112.400 ;
        RECT 148.400 112.300 149.800 112.400 ;
        RECT 146.800 111.800 149.800 112.300 ;
        RECT 150.400 111.800 151.400 112.400 ;
        RECT 157.400 112.400 158.200 119.800 ;
        RECT 158.800 113.600 159.600 114.400 ;
        RECT 159.000 112.400 159.600 113.600 ;
        RECT 157.400 111.800 158.400 112.400 ;
        RECT 159.000 112.300 160.400 112.400 ;
        RECT 161.200 112.300 162.000 119.800 ;
        RECT 159.000 111.800 162.000 112.300 ;
        RECT 165.000 118.400 165.800 119.800 ;
        RECT 165.000 117.600 166.800 118.400 ;
        RECT 165.000 112.600 165.800 117.600 ;
        RECT 170.800 115.600 171.600 119.800 ;
        RECT 174.000 115.800 174.800 119.800 ;
        RECT 174.000 115.600 174.600 115.800 ;
        RECT 171.000 115.000 174.600 115.600 ;
        RECT 172.400 112.800 173.200 114.400 ;
        RECT 165.000 111.800 166.800 112.600 ;
        RECT 174.000 112.400 174.600 115.000 ;
        RECT 175.600 113.800 176.400 119.800 ;
        RECT 175.800 113.200 176.400 113.800 ;
        RECT 178.800 119.200 182.800 119.800 ;
        RECT 178.800 113.800 179.600 119.200 ;
        RECT 180.400 113.800 181.200 118.600 ;
        RECT 182.000 114.000 182.800 119.200 ;
        RECT 183.800 119.200 187.400 119.800 ;
        RECT 183.800 119.000 184.400 119.200 ;
        RECT 178.800 113.200 179.400 113.800 ;
        RECT 175.800 112.600 179.400 113.200 ;
        RECT 180.600 113.400 181.200 113.800 ;
        RECT 183.600 113.400 184.400 119.000 ;
        RECT 186.800 119.000 187.400 119.200 ;
        RECT 180.600 113.000 184.400 113.400 ;
        RECT 185.200 113.000 186.000 118.600 ;
        RECT 186.800 113.000 187.600 119.000 ;
        RECT 180.600 112.800 184.200 113.000 ;
        RECT 185.200 112.400 185.800 113.000 ;
        RECT 188.400 112.400 189.200 119.800 ;
        RECT 146.800 111.700 149.200 111.800 ;
        RECT 146.800 111.600 147.600 111.700 ;
        RECT 148.400 111.600 149.200 111.700 ;
        RECT 138.600 110.600 142.800 111.200 ;
        RECT 138.600 110.400 139.400 110.600 ;
        RECT 140.200 109.800 141.000 110.000 ;
        RECT 137.200 109.200 141.000 109.800 ;
        RECT 137.200 109.000 138.000 109.200 ;
        RECT 107.000 107.800 118.000 108.400 ;
        RECT 107.400 107.600 108.200 107.800 ;
        RECT 110.000 107.600 110.800 107.800 ;
        RECT 100.400 106.600 104.200 107.200 ;
        RECT 98.800 104.800 99.600 106.400 ;
        RECT 100.400 102.200 101.200 106.600 ;
        RECT 103.400 106.400 104.200 106.600 ;
        RECT 113.200 105.600 113.800 107.800 ;
        RECT 116.400 107.600 118.000 107.800 ;
        RECT 121.200 107.600 122.000 108.400 ;
        RECT 125.200 107.800 136.200 108.400 ;
        RECT 125.200 107.600 126.800 107.800 ;
        RECT 111.400 105.400 112.200 105.600 ;
        RECT 105.200 104.200 106.000 105.000 ;
        RECT 109.400 104.800 112.200 105.400 ;
        RECT 113.200 104.800 114.000 105.600 ;
        RECT 109.400 104.200 110.000 104.800 ;
        RECT 114.800 104.200 115.600 105.000 ;
        RECT 104.600 103.600 106.000 104.200 ;
        RECT 104.600 102.200 105.800 103.600 ;
        RECT 109.200 102.200 110.000 104.200 ;
        RECT 113.600 103.600 115.600 104.200 ;
        RECT 113.600 102.200 114.400 103.600 ;
        RECT 118.000 102.200 118.800 107.000 ;
        RECT 121.200 104.400 121.800 107.600 ;
        RECT 122.800 104.800 123.600 106.400 ;
        RECT 121.200 102.200 122.000 104.400 ;
        RECT 124.400 102.200 125.200 107.000 ;
        RECT 129.400 105.600 130.000 107.800 ;
        RECT 135.000 107.600 135.800 107.800 ;
        RECT 142.000 107.200 142.800 110.600 ;
        RECT 150.400 108.400 151.000 111.800 ;
        RECT 151.600 110.300 152.400 110.400 ;
        RECT 156.400 110.300 157.200 110.400 ;
        RECT 151.600 109.700 157.200 110.300 ;
        RECT 151.600 108.800 152.400 109.700 ;
        RECT 156.400 108.800 157.200 109.700 ;
        RECT 157.800 110.300 158.400 111.800 ;
        RECT 159.600 111.700 162.000 111.800 ;
        RECT 159.600 111.600 160.400 111.700 ;
        RECT 159.600 110.300 160.400 110.400 ;
        RECT 157.800 109.700 160.400 110.300 ;
        RECT 157.800 108.400 158.400 109.700 ;
        RECT 159.600 109.600 160.400 109.700 ;
        RECT 148.400 107.600 151.000 108.400 ;
        RECT 153.200 108.300 154.000 108.400 ;
        RECT 154.800 108.300 155.600 108.400 ;
        RECT 153.200 108.200 155.600 108.300 ;
        RECT 152.400 107.700 156.400 108.200 ;
        RECT 152.400 107.600 154.000 107.700 ;
        RECT 154.800 107.600 156.400 107.700 ;
        RECT 157.800 107.600 160.400 108.400 ;
        RECT 139.000 106.600 142.800 107.200 ;
        RECT 139.000 106.400 139.800 106.600 ;
        RECT 127.600 104.200 128.400 105.000 ;
        RECT 129.200 104.800 130.000 105.600 ;
        RECT 131.000 105.400 131.800 105.600 ;
        RECT 131.000 104.800 133.800 105.400 ;
        RECT 133.200 104.200 133.800 104.800 ;
        RECT 137.200 104.200 138.000 105.000 ;
        RECT 142.000 104.300 142.800 106.600 ;
        RECT 143.600 106.300 144.400 106.400 ;
        RECT 148.600 106.300 149.200 107.600 ;
        RECT 152.400 107.200 153.200 107.600 ;
        RECT 155.600 107.200 156.400 107.600 ;
        RECT 143.600 105.700 149.200 106.300 ;
        RECT 150.200 106.200 153.800 106.600 ;
        RECT 155.000 106.200 158.600 106.600 ;
        RECT 159.600 106.200 160.200 107.600 ;
        RECT 143.600 105.600 144.400 105.700 ;
        RECT 145.200 104.300 146.000 104.400 ;
        RECT 127.600 103.600 129.600 104.200 ;
        RECT 128.800 102.200 129.600 103.600 ;
        RECT 133.200 102.200 134.000 104.200 ;
        RECT 137.200 103.600 138.600 104.200 ;
        RECT 137.400 102.200 138.600 103.600 ;
        RECT 142.000 103.700 146.000 104.300 ;
        RECT 142.000 102.200 142.800 103.700 ;
        RECT 145.200 103.600 146.000 103.700 ;
        RECT 148.400 102.200 149.200 105.700 ;
        RECT 150.000 106.000 154.000 106.200 ;
        RECT 150.000 102.200 150.800 106.000 ;
        RECT 153.200 102.200 154.000 106.000 ;
        RECT 154.800 106.000 158.800 106.200 ;
        RECT 154.800 102.200 155.600 106.000 ;
        RECT 158.000 102.200 158.800 106.000 ;
        RECT 159.600 102.200 160.400 106.200 ;
        RECT 161.200 102.200 162.000 111.700 ;
        RECT 164.400 109.600 165.200 111.200 ;
        RECT 166.000 108.400 166.600 111.800 ;
        RECT 169.200 110.800 170.000 112.400 ;
        RECT 174.000 111.600 174.800 112.400 ;
        RECT 185.200 112.200 186.000 112.400 ;
        RECT 182.600 111.600 186.000 112.200 ;
        RECT 188.400 111.800 190.600 112.400 ;
        RECT 170.800 109.600 172.400 110.400 ;
        RECT 174.000 108.400 174.600 111.600 ;
        RECT 180.400 109.600 182.000 110.400 ;
        RECT 166.000 107.600 166.800 108.400 ;
        RECT 173.000 108.200 174.600 108.400 ;
        RECT 172.800 107.800 174.600 108.200 ;
        RECT 175.600 108.300 176.400 108.400 ;
        RECT 178.800 108.300 180.400 108.400 ;
        RECT 162.800 106.300 163.600 106.400 ;
        RECT 164.400 106.300 165.200 106.400 ;
        RECT 162.800 105.700 165.200 106.300 ;
        RECT 162.800 104.800 163.600 105.700 ;
        RECT 164.400 105.600 165.200 105.700 ;
        RECT 166.000 104.200 166.600 107.600 ;
        RECT 167.600 104.800 168.400 106.400 ;
        RECT 166.000 102.200 166.800 104.200 ;
        RECT 172.800 102.200 173.600 107.800 ;
        RECT 175.600 107.700 180.400 108.300 ;
        RECT 175.600 107.600 176.400 107.700 ;
        RECT 178.800 107.600 180.400 107.700 ;
        RECT 182.600 105.000 183.200 111.600 ;
        RECT 190.000 111.200 190.600 111.800 ;
        RECT 190.000 110.400 191.200 111.200 ;
        RECT 188.400 108.800 189.200 110.400 ;
        RECT 190.000 107.400 190.600 110.400 ;
        RECT 179.200 104.400 183.200 105.000 ;
        RECT 179.200 104.200 179.800 104.400 ;
        RECT 178.800 103.600 179.800 104.200 ;
        RECT 182.000 104.200 183.200 104.400 ;
        RECT 188.400 106.800 190.600 107.400 ;
        RECT 178.800 102.200 179.600 103.600 ;
        RECT 182.000 102.200 182.800 104.200 ;
        RECT 188.400 102.200 189.200 106.800 ;
        RECT 4.400 95.200 5.200 99.800 ;
        RECT 3.000 94.600 5.200 95.200 ;
        RECT 6.000 95.400 6.800 99.800 ;
        RECT 10.200 98.400 11.400 99.800 ;
        RECT 10.200 97.800 11.600 98.400 ;
        RECT 14.800 97.800 15.600 99.800 ;
        RECT 19.200 98.400 20.000 99.800 ;
        RECT 19.200 97.800 21.200 98.400 ;
        RECT 10.800 97.000 11.600 97.800 ;
        RECT 15.000 97.200 15.600 97.800 ;
        RECT 15.000 96.600 17.800 97.200 ;
        RECT 17.000 96.400 17.800 96.600 ;
        RECT 18.800 96.400 19.600 97.200 ;
        RECT 20.400 97.000 21.200 97.800 ;
        RECT 12.400 96.300 13.200 96.400 ;
        RECT 9.200 95.700 13.200 96.300 ;
        RECT 9.200 95.600 10.000 95.700 ;
        RECT 12.400 95.600 13.200 95.700 ;
        RECT 9.000 95.400 10.000 95.600 ;
        RECT 6.000 94.800 10.000 95.400 ;
        RECT 3.000 91.600 3.600 94.600 ;
        RECT 4.400 92.300 5.200 93.200 ;
        RECT 6.000 92.300 6.800 94.800 ;
        RECT 13.000 94.200 13.800 94.400 ;
        RECT 17.200 94.200 18.000 94.400 ;
        RECT 18.800 94.200 19.400 96.400 ;
        RECT 23.600 95.000 24.400 99.800 ;
        RECT 25.200 96.000 26.000 99.800 ;
        RECT 28.400 96.000 29.200 99.800 ;
        RECT 25.200 95.800 29.200 96.000 ;
        RECT 30.000 95.800 30.800 99.800 ;
        RECT 33.200 97.800 34.000 99.800 ;
        RECT 25.400 95.400 29.000 95.800 ;
        RECT 26.000 94.400 26.800 94.800 ;
        RECT 30.000 94.400 30.600 95.800 ;
        RECT 33.200 94.400 33.800 97.800 ;
        RECT 38.000 97.600 38.800 99.800 ;
        RECT 34.800 96.300 35.600 97.200 ;
        RECT 38.000 96.300 38.600 97.600 ;
        RECT 34.800 95.700 38.700 96.300 ;
        RECT 34.800 95.600 35.600 95.700 ;
        RECT 38.000 94.400 38.600 95.700 ;
        RECT 39.600 95.600 40.400 97.200 ;
        RECT 41.200 95.600 42.000 97.200 ;
        RECT 22.000 94.200 23.600 94.400 ;
        RECT 12.600 93.600 23.600 94.200 ;
        RECT 25.200 93.800 26.800 94.400 ;
        RECT 25.200 93.600 26.000 93.800 ;
        RECT 28.200 93.600 30.800 94.400 ;
        RECT 31.600 94.300 32.400 94.400 ;
        RECT 33.200 94.300 34.000 94.400 ;
        RECT 31.600 93.700 34.000 94.300 ;
        RECT 31.600 93.600 32.400 93.700 ;
        RECT 33.200 93.600 34.000 93.700 ;
        RECT 38.000 93.600 38.800 94.400 ;
        RECT 42.800 94.300 43.600 99.800 ;
        RECT 47.000 98.400 47.800 99.800 ;
        RECT 46.000 97.600 47.800 98.400 ;
        RECT 47.000 96.400 47.800 97.600 ;
        RECT 46.000 95.800 47.800 96.400 ;
        RECT 44.400 94.300 45.200 95.200 ;
        RECT 42.800 93.700 45.200 94.300 ;
        RECT 10.800 92.800 11.600 93.000 ;
        RECT 4.400 91.700 6.800 92.300 ;
        RECT 7.800 92.200 11.600 92.800 ;
        RECT 7.800 92.000 8.600 92.200 ;
        RECT 4.400 91.600 5.200 91.700 ;
        RECT 2.400 90.800 3.600 91.600 ;
        RECT 3.000 90.200 3.600 90.800 ;
        RECT 6.000 91.400 6.800 91.700 ;
        RECT 9.400 91.400 10.200 91.600 ;
        RECT 6.000 90.800 10.200 91.400 ;
        RECT 3.000 89.600 5.200 90.200 ;
        RECT 4.400 82.200 5.200 89.600 ;
        RECT 6.000 82.200 6.800 90.800 ;
        RECT 12.600 90.400 13.200 93.600 ;
        RECT 19.800 93.400 20.600 93.600 ;
        RECT 18.800 92.400 19.600 92.600 ;
        RECT 21.400 92.400 22.200 92.600 ;
        RECT 17.200 91.800 22.200 92.400 ;
        RECT 17.200 91.600 18.000 91.800 ;
        RECT 26.800 91.600 27.600 93.200 ;
        RECT 28.200 92.300 28.800 93.600 ;
        RECT 31.600 92.300 32.400 92.400 ;
        RECT 28.200 91.700 32.400 92.300 ;
        RECT 18.800 91.000 24.400 91.200 ;
        RECT 18.600 90.800 24.400 91.000 ;
        RECT 10.800 89.800 13.200 90.400 ;
        RECT 14.600 90.600 24.400 90.800 ;
        RECT 14.600 90.200 19.400 90.600 ;
        RECT 10.800 88.800 11.400 89.800 ;
        RECT 10.000 88.000 11.400 88.800 ;
        RECT 13.000 89.000 13.800 89.200 ;
        RECT 14.600 89.000 15.200 90.200 ;
        RECT 13.000 88.400 15.200 89.000 ;
        RECT 15.800 89.000 21.200 89.600 ;
        RECT 15.800 88.800 16.600 89.000 ;
        RECT 20.400 88.800 21.200 89.000 ;
        RECT 14.200 87.400 15.000 87.600 ;
        RECT 17.000 87.400 17.800 87.600 ;
        RECT 10.800 86.200 11.600 87.000 ;
        RECT 14.200 86.800 17.800 87.400 ;
        RECT 15.000 86.200 15.600 86.800 ;
        RECT 20.400 86.200 21.200 87.000 ;
        RECT 10.200 82.200 11.400 86.200 ;
        RECT 14.800 82.200 15.600 86.200 ;
        RECT 19.200 85.600 21.200 86.200 ;
        RECT 19.200 82.200 20.000 85.600 ;
        RECT 23.600 82.200 24.400 90.600 ;
        RECT 28.200 90.200 28.800 91.700 ;
        RECT 31.600 90.800 32.400 91.700 ;
        RECT 30.000 90.200 30.800 90.400 ;
        RECT 33.200 90.200 33.800 93.600 ;
        RECT 36.400 90.800 37.200 92.400 ;
        RECT 38.000 90.200 38.600 93.600 ;
        RECT 42.800 92.300 43.600 93.700 ;
        RECT 44.400 93.600 45.200 93.700 ;
        RECT 44.400 92.300 45.200 92.400 ;
        RECT 42.800 91.700 45.200 92.300 ;
        RECT 27.800 89.600 28.800 90.200 ;
        RECT 29.400 89.600 30.800 90.200 ;
        RECT 27.800 82.200 28.600 89.600 ;
        RECT 29.400 88.400 30.000 89.600 ;
        RECT 29.200 87.600 30.000 88.400 ;
        RECT 32.200 89.400 34.000 90.200 ;
        RECT 37.000 89.400 38.800 90.200 ;
        RECT 32.200 82.200 33.000 89.400 ;
        RECT 37.000 82.200 37.800 89.400 ;
        RECT 42.800 82.200 43.600 91.700 ;
        RECT 44.400 91.600 45.200 91.700 ;
        RECT 46.000 82.200 46.800 95.800 ;
        RECT 49.200 92.400 50.000 99.800 ;
        RECT 52.400 95.200 53.200 99.800 ;
        RECT 58.800 95.800 59.600 99.800 ;
        RECT 63.000 98.400 63.800 99.800 ;
        RECT 63.000 97.600 64.400 98.400 ;
        RECT 63.000 96.800 63.800 97.600 ;
        RECT 63.000 95.800 64.400 96.800 ;
        RECT 67.800 96.400 68.600 99.800 ;
        RECT 51.000 94.600 53.200 95.200 ;
        RECT 59.000 95.600 59.600 95.800 ;
        RECT 59.000 95.200 60.800 95.600 ;
        RECT 59.000 95.000 63.200 95.200 ;
        RECT 60.200 94.600 63.200 95.000 ;
        RECT 47.600 88.800 48.400 90.400 ;
        RECT 49.200 90.200 49.800 92.400 ;
        RECT 51.000 91.600 51.600 94.600 ;
        RECT 62.400 94.400 63.200 94.600 ;
        RECT 52.400 92.300 53.200 93.200 ;
        RECT 58.800 92.800 59.600 94.400 ;
        RECT 60.800 93.800 61.600 94.000 ;
        RECT 60.600 93.200 61.600 93.800 ;
        RECT 60.600 92.400 61.200 93.200 ;
        RECT 54.000 92.300 54.800 92.400 ;
        RECT 52.400 91.700 54.800 92.300 ;
        RECT 52.400 91.600 53.200 91.700 ;
        RECT 54.000 91.600 54.800 91.700 ;
        RECT 60.400 91.600 61.200 92.400 ;
        RECT 50.400 90.800 51.600 91.600 ;
        RECT 62.400 91.000 63.000 94.400 ;
        RECT 63.800 92.400 64.400 95.800 ;
        RECT 63.600 91.600 64.400 92.400 ;
        RECT 51.000 90.200 51.600 90.800 ;
        RECT 60.600 90.400 63.000 91.000 ;
        RECT 49.200 82.200 50.000 90.200 ;
        RECT 51.000 89.600 53.200 90.200 ;
        RECT 52.400 82.200 53.200 89.600 ;
        RECT 60.600 86.200 61.200 90.400 ;
        RECT 63.800 90.200 64.400 91.600 ;
        RECT 60.400 82.200 61.200 86.200 ;
        RECT 63.600 82.200 64.400 90.200 ;
        RECT 66.800 95.800 68.600 96.400 ;
        RECT 71.600 97.800 72.400 99.800 ;
        RECT 66.800 92.300 67.600 95.800 ;
        RECT 71.600 94.400 72.200 97.800 ;
        RECT 73.200 95.600 74.000 97.200 ;
        RECT 70.000 94.300 70.800 94.400 ;
        RECT 71.600 94.300 72.400 94.400 ;
        RECT 70.000 93.700 72.400 94.300 ;
        RECT 70.000 93.600 70.800 93.700 ;
        RECT 71.600 93.600 72.400 93.700 ;
        RECT 70.000 92.300 70.800 92.400 ;
        RECT 66.800 91.700 70.800 92.300 ;
        RECT 66.800 82.200 67.600 91.700 ;
        RECT 70.000 90.800 70.800 91.700 ;
        RECT 68.400 88.800 69.200 90.400 ;
        RECT 71.600 90.200 72.200 93.600 ;
        RECT 74.800 92.400 75.600 99.800 ;
        RECT 78.000 95.200 78.800 99.800 ;
        RECT 76.600 94.600 78.800 95.200 ;
        RECT 81.200 97.800 82.000 99.800 ;
        RECT 86.000 97.800 86.800 99.800 ;
        RECT 74.800 90.200 75.400 92.400 ;
        RECT 76.600 91.600 77.200 94.600 ;
        RECT 81.200 94.400 81.800 97.800 ;
        RECT 82.800 96.300 83.600 97.200 ;
        RECT 84.400 96.300 85.200 96.400 ;
        RECT 82.800 95.700 85.200 96.300 ;
        RECT 82.800 95.600 83.600 95.700 ;
        RECT 84.400 95.600 85.200 95.700 ;
        RECT 86.000 94.400 86.600 97.800 ;
        RECT 87.600 95.600 88.400 97.200 ;
        RECT 89.200 95.400 90.000 99.800 ;
        RECT 93.400 98.400 94.600 99.800 ;
        RECT 93.400 97.800 94.800 98.400 ;
        RECT 98.000 97.800 98.800 99.800 ;
        RECT 102.400 98.400 103.200 99.800 ;
        RECT 102.400 97.800 104.400 98.400 ;
        RECT 94.000 97.000 94.800 97.800 ;
        RECT 98.200 97.200 98.800 97.800 ;
        RECT 98.200 96.600 101.000 97.200 ;
        RECT 100.200 96.400 101.000 96.600 ;
        RECT 102.000 96.400 102.800 97.200 ;
        RECT 103.600 97.000 104.400 97.800 ;
        RECT 92.200 95.400 93.000 95.600 ;
        RECT 89.200 94.800 93.000 95.400 ;
        RECT 81.200 93.600 82.000 94.400 ;
        RECT 86.000 93.600 86.800 94.400 ;
        RECT 78.000 91.600 78.800 93.200 ;
        RECT 76.000 90.800 77.200 91.600 ;
        RECT 79.600 90.800 80.400 92.400 ;
        RECT 81.200 92.300 81.800 93.600 ;
        RECT 84.400 92.300 85.200 92.400 ;
        RECT 81.200 91.700 85.200 92.300 ;
        RECT 76.600 90.200 77.200 90.800 ;
        RECT 81.200 90.200 81.800 91.700 ;
        RECT 84.400 90.800 85.200 91.700 ;
        RECT 86.000 92.300 86.600 93.600 ;
        RECT 87.600 92.300 88.400 92.400 ;
        RECT 86.000 91.700 88.400 92.300 ;
        RECT 86.000 90.200 86.600 91.700 ;
        RECT 87.600 91.600 88.400 91.700 ;
        RECT 89.200 91.400 90.000 94.800 ;
        RECT 96.200 94.200 97.000 94.400 ;
        RECT 102.000 94.200 102.600 96.400 ;
        RECT 106.800 95.000 107.600 99.800 ;
        RECT 108.400 95.200 109.200 99.800 ;
        RECT 108.400 94.600 110.600 95.200 ;
        RECT 105.200 94.200 106.800 94.400 ;
        RECT 95.800 93.600 106.800 94.200 ;
        RECT 94.000 92.800 94.800 93.000 ;
        RECT 91.000 92.200 94.800 92.800 ;
        RECT 95.800 92.400 96.400 93.600 ;
        RECT 103.000 93.400 103.800 93.600 ;
        RECT 104.600 92.400 105.400 92.600 ;
        RECT 91.000 92.000 91.800 92.200 ;
        RECT 95.600 91.600 96.400 92.400 ;
        RECT 98.800 92.300 99.600 92.400 ;
        RECT 100.400 92.300 105.400 92.400 ;
        RECT 98.800 91.800 105.400 92.300 ;
        RECT 98.800 91.700 101.200 91.800 ;
        RECT 98.800 91.600 99.600 91.700 ;
        RECT 100.400 91.600 101.200 91.700 ;
        RECT 108.400 91.600 109.200 93.200 ;
        RECT 110.000 91.600 110.600 94.600 ;
        RECT 111.600 92.400 112.400 99.800 ;
        RECT 92.600 91.400 93.400 91.600 ;
        RECT 89.200 90.800 93.400 91.400 ;
        RECT 70.600 89.400 72.400 90.200 ;
        RECT 70.600 82.200 71.400 89.400 ;
        RECT 74.800 82.200 75.600 90.200 ;
        RECT 76.600 89.600 78.800 90.200 ;
        RECT 78.000 82.200 78.800 89.600 ;
        RECT 80.200 89.400 82.000 90.200 ;
        RECT 85.000 89.400 86.800 90.200 ;
        RECT 80.200 82.200 81.000 89.400 ;
        RECT 85.000 82.200 85.800 89.400 ;
        RECT 89.200 82.200 90.000 90.800 ;
        RECT 95.800 90.400 96.400 91.600 ;
        RECT 102.000 91.000 107.600 91.200 ;
        RECT 101.800 90.800 107.600 91.000 ;
        RECT 94.000 89.800 96.400 90.400 ;
        RECT 97.800 90.600 107.600 90.800 ;
        RECT 97.800 90.200 102.600 90.600 ;
        RECT 94.000 88.800 94.600 89.800 ;
        RECT 93.200 88.000 94.600 88.800 ;
        RECT 96.200 89.000 97.000 89.200 ;
        RECT 97.800 89.000 98.400 90.200 ;
        RECT 96.200 88.400 98.400 89.000 ;
        RECT 99.000 89.000 104.400 89.600 ;
        RECT 99.000 88.800 99.800 89.000 ;
        RECT 103.600 88.800 104.400 89.000 ;
        RECT 97.400 87.400 98.200 87.600 ;
        RECT 100.200 87.400 101.000 87.600 ;
        RECT 94.000 86.200 94.800 87.000 ;
        RECT 97.400 86.800 101.000 87.400 ;
        RECT 98.200 86.200 98.800 86.800 ;
        RECT 103.600 86.200 104.400 87.000 ;
        RECT 93.400 82.200 94.600 86.200 ;
        RECT 98.000 82.200 98.800 86.200 ;
        RECT 102.400 85.600 104.400 86.200 ;
        RECT 102.400 82.200 103.200 85.600 ;
        RECT 106.800 82.200 107.600 90.600 ;
        RECT 110.000 90.800 111.200 91.600 ;
        RECT 110.000 90.200 110.600 90.800 ;
        RECT 111.800 90.200 112.400 92.400 ;
        RECT 108.400 89.600 110.600 90.200 ;
        RECT 108.400 82.200 109.200 89.600 ;
        RECT 111.600 82.200 112.400 90.200 ;
        RECT 113.200 94.300 114.000 99.800 ;
        RECT 114.800 95.600 115.600 97.200 ;
        RECT 114.800 94.300 115.600 94.400 ;
        RECT 113.200 93.700 115.600 94.300 ;
        RECT 113.200 82.200 114.000 93.700 ;
        RECT 114.800 93.600 115.600 93.700 ;
        RECT 114.800 88.300 115.600 88.400 ;
        RECT 116.400 88.300 117.200 99.800 ;
        RECT 118.000 95.600 118.800 97.200 ;
        RECT 122.800 95.800 123.600 99.800 ;
        RECT 124.200 96.400 125.000 97.200 ;
        RECT 121.200 92.800 122.000 94.400 ;
        RECT 119.600 92.200 120.400 92.400 ;
        RECT 122.800 92.200 123.400 95.800 ;
        RECT 124.400 95.600 125.200 96.400 ;
        RECT 127.200 94.200 128.000 99.800 ;
        RECT 135.600 95.800 136.400 99.800 ;
        RECT 137.000 96.400 137.800 97.200 ;
        RECT 126.200 93.800 128.000 94.200 ;
        RECT 126.200 93.600 127.800 93.800 ;
        RECT 126.200 92.400 126.800 93.600 ;
        RECT 134.000 92.800 134.800 94.400 ;
        RECT 135.600 94.300 136.200 95.800 ;
        RECT 137.200 95.600 138.000 96.400 ;
        RECT 143.600 95.600 144.400 97.200 ;
        RECT 142.000 94.300 142.800 94.400 ;
        RECT 135.600 93.700 142.800 94.300 ;
        RECT 124.400 92.200 125.200 92.400 ;
        RECT 119.600 91.600 121.200 92.200 ;
        RECT 122.800 91.600 125.200 92.200 ;
        RECT 126.000 91.600 126.800 92.400 ;
        RECT 128.400 91.600 130.000 92.400 ;
        RECT 120.400 91.200 121.200 91.600 ;
        RECT 124.400 90.200 125.000 91.600 ;
        RECT 126.200 90.400 126.800 91.600 ;
        RECT 114.800 87.700 117.200 88.300 ;
        RECT 114.800 87.600 115.600 87.700 ;
        RECT 116.400 82.200 117.200 87.700 ;
        RECT 119.600 89.600 123.600 90.200 ;
        RECT 119.600 82.200 120.400 89.600 ;
        RECT 122.800 82.200 123.600 89.600 ;
        RECT 124.400 82.200 125.200 90.200 ;
        RECT 126.000 89.600 126.800 90.400 ;
        RECT 130.800 89.600 131.600 92.400 ;
        RECT 132.400 92.200 133.200 92.400 ;
        RECT 135.600 92.200 136.200 93.700 ;
        RECT 142.000 93.600 142.800 93.700 ;
        RECT 137.200 92.200 138.000 92.400 ;
        RECT 132.400 91.600 134.000 92.200 ;
        RECT 135.600 91.600 138.000 92.200 ;
        RECT 133.200 91.200 134.000 91.600 ;
        RECT 137.200 90.200 137.800 91.600 ;
        RECT 132.400 89.600 136.400 90.200 ;
        RECT 126.200 87.000 126.800 89.600 ;
        RECT 127.600 87.600 128.400 89.200 ;
        RECT 126.200 86.400 129.800 87.000 ;
        RECT 126.200 86.200 126.800 86.400 ;
        RECT 126.000 82.200 126.800 86.200 ;
        RECT 129.200 86.200 129.800 86.400 ;
        RECT 129.200 82.200 130.000 86.200 ;
        RECT 132.400 82.200 133.200 89.600 ;
        RECT 135.600 82.200 136.400 89.600 ;
        RECT 137.200 82.200 138.000 90.200 ;
        RECT 145.200 82.200 146.000 99.800 ;
        RECT 146.800 95.800 147.600 99.800 ;
        RECT 148.400 96.000 149.200 99.800 ;
        RECT 151.600 96.000 152.400 99.800 ;
        RECT 153.400 96.400 154.200 97.200 ;
        RECT 148.400 95.800 152.400 96.000 ;
        RECT 147.000 94.400 147.600 95.800 ;
        RECT 148.600 95.400 152.200 95.800 ;
        RECT 153.200 95.600 154.000 96.400 ;
        RECT 154.800 95.800 155.600 99.800 ;
        RECT 150.800 94.400 151.600 94.800 ;
        RECT 146.800 93.600 149.400 94.400 ;
        RECT 150.800 93.800 152.400 94.400 ;
        RECT 151.600 93.600 152.400 93.800 ;
        RECT 146.800 90.200 147.600 90.400 ;
        RECT 148.800 90.200 149.400 93.600 ;
        RECT 150.000 91.600 150.800 93.200 ;
        RECT 153.200 92.200 154.000 92.400 ;
        RECT 155.000 92.200 155.600 95.800 ;
        RECT 159.600 95.600 160.400 97.200 ;
        RECT 161.200 96.300 162.000 99.800 ;
        RECT 166.000 98.400 166.800 99.800 ;
        RECT 166.000 97.800 167.000 98.400 ;
        RECT 166.400 97.600 167.000 97.800 ;
        RECT 169.200 98.300 170.000 99.800 ;
        RECT 174.000 98.300 174.800 98.400 ;
        RECT 169.200 97.700 174.800 98.300 ;
        RECT 169.200 97.600 170.400 97.700 ;
        RECT 174.000 97.600 174.800 97.700 ;
        RECT 166.400 97.000 170.400 97.600 ;
        RECT 164.400 96.300 166.200 96.400 ;
        RECT 161.200 95.700 166.200 96.300 ;
        RECT 156.400 92.800 157.200 94.400 ;
        RECT 158.000 92.200 158.800 92.400 ;
        RECT 153.200 91.600 155.600 92.200 ;
        RECT 157.200 91.600 158.800 92.200 ;
        RECT 153.400 90.200 154.000 91.600 ;
        RECT 157.200 91.200 158.000 91.600 ;
        RECT 146.800 89.600 148.200 90.200 ;
        RECT 148.800 89.600 149.800 90.200 ;
        RECT 147.600 88.400 148.200 89.600 ;
        RECT 147.600 87.600 148.400 88.400 ;
        RECT 149.000 82.200 149.800 89.600 ;
        RECT 153.200 82.200 154.000 90.200 ;
        RECT 154.800 89.600 158.800 90.200 ;
        RECT 154.800 82.200 155.600 89.600 ;
        RECT 158.000 82.200 158.800 89.600 ;
        RECT 161.200 82.200 162.000 95.700 ;
        RECT 164.400 95.600 166.200 95.700 ;
        RECT 166.000 93.600 167.600 94.400 ;
        RECT 164.400 92.300 165.200 92.400 ;
        RECT 167.600 92.300 169.200 92.400 ;
        RECT 164.400 91.700 169.200 92.300 ;
        RECT 164.400 91.600 165.200 91.700 ;
        RECT 167.600 91.600 169.200 91.700 ;
        RECT 169.800 90.400 170.400 97.000 ;
        RECT 175.600 95.200 176.400 99.800 ;
        RECT 175.600 94.600 177.800 95.200 ;
        RECT 172.400 92.300 173.200 92.400 ;
        RECT 175.600 92.300 176.400 93.200 ;
        RECT 172.400 91.700 176.400 92.300 ;
        RECT 172.400 91.600 173.200 91.700 ;
        RECT 175.600 91.600 176.400 91.700 ;
        RECT 177.200 91.600 177.800 94.600 ;
        RECT 177.200 90.800 178.400 91.600 ;
        RECT 169.800 89.800 173.200 90.400 ;
        RECT 177.200 90.200 177.800 90.800 ;
        RECT 172.400 89.600 173.200 89.800 ;
        RECT 175.600 89.600 177.800 90.200 ;
        RECT 163.000 88.800 166.600 89.400 ;
        RECT 163.000 88.200 163.600 88.800 ;
        RECT 162.800 82.200 163.600 88.200 ;
        RECT 166.000 88.200 166.600 88.800 ;
        RECT 167.800 89.000 171.400 89.200 ;
        RECT 172.400 89.000 173.000 89.600 ;
        RECT 167.800 88.600 171.600 89.000 ;
        RECT 167.800 88.200 168.400 88.600 ;
        RECT 166.000 82.800 166.800 88.200 ;
        RECT 167.600 83.400 168.400 88.200 ;
        RECT 169.200 82.800 170.000 88.000 ;
        RECT 170.800 83.000 171.600 88.600 ;
        RECT 172.400 83.400 173.200 89.000 ;
        RECT 166.000 82.200 170.000 82.800 ;
        RECT 171.000 82.800 171.600 83.000 ;
        RECT 174.000 83.000 174.800 89.000 ;
        RECT 174.000 82.800 174.600 83.000 ;
        RECT 171.000 82.200 174.600 82.800 ;
        RECT 175.600 82.200 176.400 89.600 ;
        RECT 180.400 82.200 181.200 99.800 ;
        RECT 182.000 95.600 182.800 97.200 ;
        RECT 183.600 95.200 184.400 99.800 ;
        RECT 188.400 95.200 189.200 99.800 ;
        RECT 183.600 94.600 185.800 95.200 ;
        RECT 188.400 94.600 190.600 95.200 ;
        RECT 183.600 91.600 184.400 93.200 ;
        RECT 185.200 91.600 185.800 94.600 ;
        RECT 188.400 91.600 189.200 93.200 ;
        RECT 190.000 91.600 190.600 94.600 ;
        RECT 185.200 90.800 186.400 91.600 ;
        RECT 190.000 90.800 191.200 91.600 ;
        RECT 185.200 90.200 185.800 90.800 ;
        RECT 190.000 90.200 190.600 90.800 ;
        RECT 183.600 89.600 185.800 90.200 ;
        RECT 188.400 89.600 190.600 90.200 ;
        RECT 183.600 82.200 184.400 89.600 ;
        RECT 188.400 82.200 189.200 89.600 ;
        RECT 4.400 72.400 5.200 79.800 ;
        RECT 6.000 75.800 6.800 79.800 ;
        RECT 6.200 75.600 6.800 75.800 ;
        RECT 9.200 75.800 10.000 79.800 ;
        RECT 9.200 75.600 9.800 75.800 ;
        RECT 6.200 75.000 9.800 75.600 ;
        RECT 6.200 72.400 6.800 75.000 ;
        RECT 7.600 72.800 8.400 74.400 ;
        RECT 15.000 72.400 15.800 79.800 ;
        RECT 16.400 73.600 17.200 74.400 ;
        RECT 16.600 72.400 17.200 73.600 ;
        RECT 19.400 72.600 20.200 79.800 ;
        RECT 3.000 71.800 5.200 72.400 ;
        RECT 3.000 71.200 3.600 71.800 ;
        RECT 6.000 71.600 6.800 72.400 ;
        RECT 2.400 70.400 3.600 71.200 ;
        RECT 3.000 67.400 3.600 70.400 ;
        RECT 4.400 68.800 5.200 70.400 ;
        RECT 6.200 68.400 6.800 71.600 ;
        RECT 10.800 70.800 11.600 72.400 ;
        RECT 15.000 71.800 16.000 72.400 ;
        RECT 16.600 71.800 18.000 72.400 ;
        RECT 19.400 71.800 21.200 72.600 ;
        RECT 8.400 69.600 10.000 70.400 ;
        RECT 14.000 68.800 14.800 70.400 ;
        RECT 15.400 70.300 16.000 71.800 ;
        RECT 17.200 71.600 18.000 71.800 ;
        RECT 18.800 70.300 19.600 71.200 ;
        RECT 15.400 69.700 19.600 70.300 ;
        RECT 15.400 68.400 16.000 69.700 ;
        RECT 18.800 69.600 19.600 69.700 ;
        RECT 20.400 68.400 21.000 71.800 ;
        RECT 6.200 68.200 7.800 68.400 ;
        RECT 6.200 67.800 8.000 68.200 ;
        RECT 3.000 66.800 5.200 67.400 ;
        RECT 4.400 62.200 5.200 66.800 ;
        RECT 7.200 62.200 8.000 67.800 ;
        RECT 15.400 67.600 18.000 68.400 ;
        RECT 20.400 67.600 21.200 68.400 ;
        RECT 12.600 66.200 16.200 66.600 ;
        RECT 17.200 66.200 17.800 67.600 ;
        RECT 18.800 66.300 19.600 66.400 ;
        RECT 20.400 66.300 21.000 67.600 ;
        RECT 23.600 66.800 24.400 68.400 ;
        RECT 12.400 66.000 16.400 66.200 ;
        RECT 12.400 62.200 13.200 66.000 ;
        RECT 15.600 62.200 16.400 66.000 ;
        RECT 17.200 62.200 18.000 66.200 ;
        RECT 18.800 65.700 21.100 66.300 ;
        RECT 18.800 65.600 19.600 65.700 ;
        RECT 20.400 64.200 21.000 65.700 ;
        RECT 22.000 64.800 22.800 66.400 ;
        RECT 25.200 66.300 26.000 79.800 ;
        RECT 26.800 71.600 27.600 73.200 ;
        RECT 28.400 66.300 29.200 66.400 ;
        RECT 25.200 65.700 29.200 66.300 ;
        RECT 25.200 65.600 27.000 65.700 ;
        RECT 20.400 62.200 21.200 64.200 ;
        RECT 26.200 62.200 27.000 65.600 ;
        RECT 28.400 64.800 29.200 65.700 ;
        RECT 30.000 62.200 30.800 79.800 ;
        RECT 34.200 72.400 35.000 79.800 ;
        RECT 35.600 73.600 36.400 74.400 ;
        RECT 35.800 72.400 36.400 73.600 ;
        RECT 38.600 72.600 39.400 79.800 ;
        RECT 34.200 71.800 35.200 72.400 ;
        RECT 35.800 71.800 37.200 72.400 ;
        RECT 38.600 71.800 40.400 72.600 ;
        RECT 33.200 68.800 34.000 70.400 ;
        RECT 34.600 68.400 35.200 71.800 ;
        RECT 36.400 71.600 37.200 71.800 ;
        RECT 39.600 71.600 40.400 71.800 ;
        RECT 38.000 69.600 38.800 71.200 ;
        RECT 39.600 68.400 40.200 71.600 ;
        RECT 42.800 71.400 43.600 79.800 ;
        RECT 47.200 76.400 48.000 79.800 ;
        RECT 46.000 75.800 48.000 76.400 ;
        RECT 51.600 75.800 52.400 79.800 ;
        RECT 55.800 75.800 57.000 79.800 ;
        RECT 46.000 75.000 46.800 75.800 ;
        RECT 51.600 75.200 52.200 75.800 ;
        RECT 49.400 74.600 53.000 75.200 ;
        RECT 55.600 75.000 56.400 75.800 ;
        RECT 49.400 74.400 50.200 74.600 ;
        RECT 52.200 74.400 53.000 74.600 ;
        RECT 46.000 73.000 46.800 73.200 ;
        RECT 50.600 73.000 51.400 73.200 ;
        RECT 46.000 72.400 51.400 73.000 ;
        RECT 52.000 73.000 54.200 73.600 ;
        RECT 52.000 71.800 52.600 73.000 ;
        RECT 53.400 72.800 54.200 73.000 ;
        RECT 55.800 73.200 57.200 74.000 ;
        RECT 55.800 72.200 56.400 73.200 ;
        RECT 47.800 71.400 52.600 71.800 ;
        RECT 42.800 71.200 52.600 71.400 ;
        RECT 54.000 71.600 56.400 72.200 ;
        RECT 42.800 71.000 48.600 71.200 ;
        RECT 42.800 70.800 48.400 71.000 ;
        RECT 49.200 70.200 50.000 70.400 ;
        RECT 45.000 69.600 50.000 70.200 ;
        RECT 45.000 69.400 45.800 69.600 ;
        RECT 47.600 69.400 48.400 69.600 ;
        RECT 46.600 68.400 47.400 68.600 ;
        RECT 54.000 68.400 54.600 71.600 ;
        RECT 60.400 71.200 61.200 79.800 ;
        RECT 57.000 70.600 61.200 71.200 ;
        RECT 57.000 70.400 57.800 70.600 ;
        RECT 58.600 69.800 59.400 70.000 ;
        RECT 55.600 69.200 59.400 69.800 ;
        RECT 55.600 69.000 56.400 69.200 ;
        RECT 31.600 68.200 32.400 68.400 ;
        RECT 31.600 67.600 33.200 68.200 ;
        RECT 34.600 67.600 37.200 68.400 ;
        RECT 39.600 67.600 40.400 68.400 ;
        RECT 43.600 67.800 54.600 68.400 ;
        RECT 43.600 67.600 45.200 67.800 ;
        RECT 32.400 67.200 33.200 67.600 ;
        RECT 31.800 66.200 35.400 66.600 ;
        RECT 36.400 66.300 37.000 67.600 ;
        RECT 38.000 66.300 38.800 66.400 ;
        RECT 31.600 66.000 35.600 66.200 ;
        RECT 31.600 62.200 32.400 66.000 ;
        RECT 34.800 62.200 35.600 66.000 ;
        RECT 36.400 65.700 38.800 66.300 ;
        RECT 36.400 62.200 37.200 65.700 ;
        RECT 38.000 65.600 38.800 65.700 ;
        RECT 39.600 64.200 40.200 67.600 ;
        RECT 41.200 64.800 42.000 66.400 ;
        RECT 39.600 62.200 40.400 64.200 ;
        RECT 42.800 62.200 43.600 67.000 ;
        RECT 47.800 66.400 48.400 67.800 ;
        RECT 53.400 67.600 54.200 67.800 ;
        RECT 60.400 67.200 61.200 70.600 ;
        RECT 57.400 66.600 61.200 67.200 ;
        RECT 57.400 66.400 58.200 66.600 ;
        RECT 46.000 64.200 46.800 65.000 ;
        RECT 47.600 64.800 48.400 66.400 ;
        RECT 49.400 65.400 50.200 65.600 ;
        RECT 49.400 64.800 52.200 65.400 ;
        RECT 51.600 64.200 52.200 64.800 ;
        RECT 55.600 64.200 56.400 65.000 ;
        RECT 46.000 63.600 48.000 64.200 ;
        RECT 47.200 62.200 48.000 63.600 ;
        RECT 51.600 62.200 52.400 64.200 ;
        RECT 55.600 63.600 57.000 64.200 ;
        RECT 55.800 62.200 57.000 63.600 ;
        RECT 60.400 62.200 61.200 66.600 ;
        RECT 68.400 62.200 69.200 79.800 ;
        RECT 70.000 71.800 70.800 79.800 ;
        RECT 73.200 72.400 74.000 79.800 ;
        RECT 71.800 71.800 74.000 72.400 ;
        RECT 70.000 69.600 70.600 71.800 ;
        RECT 71.800 71.200 72.400 71.800 ;
        RECT 71.200 70.400 72.400 71.200 ;
        RECT 76.400 71.200 77.200 79.800 ;
        RECT 79.600 71.200 80.400 79.800 ;
        RECT 82.800 71.200 83.600 79.800 ;
        RECT 86.000 71.200 86.800 79.800 ;
        RECT 89.200 72.400 90.000 79.800 ;
        RECT 92.400 74.300 93.200 79.800 ;
        RECT 94.800 74.300 95.600 74.400 ;
        RECT 92.400 73.700 95.600 74.300 ;
        RECT 89.200 71.800 91.400 72.400 ;
        RECT 92.400 71.800 93.200 73.700 ;
        RECT 94.800 73.600 95.600 73.700 ;
        RECT 94.800 72.400 95.400 73.600 ;
        RECT 96.200 72.400 97.000 79.800 ;
        RECT 90.800 71.200 91.400 71.800 ;
        RECT 76.400 70.400 78.200 71.200 ;
        RECT 79.600 70.400 81.800 71.200 ;
        RECT 82.800 70.400 85.000 71.200 ;
        RECT 86.000 70.400 88.400 71.200 ;
        RECT 90.800 70.400 92.000 71.200 ;
        RECT 70.000 62.200 70.800 69.600 ;
        RECT 71.800 67.400 72.400 70.400 ;
        RECT 73.200 68.800 74.000 70.400 ;
        RECT 77.400 69.000 78.200 70.400 ;
        RECT 81.000 69.000 81.800 70.400 ;
        RECT 84.200 69.000 85.000 70.400 ;
        RECT 77.400 68.200 80.000 69.000 ;
        RECT 81.000 68.200 83.400 69.000 ;
        RECT 84.200 68.200 86.800 69.000 ;
        RECT 77.400 67.600 78.200 68.200 ;
        RECT 81.000 67.600 81.800 68.200 ;
        RECT 84.200 67.600 85.000 68.200 ;
        RECT 87.600 67.600 88.400 70.400 ;
        RECT 89.200 68.800 90.000 70.400 ;
        RECT 71.800 66.800 74.000 67.400 ;
        RECT 73.200 62.200 74.000 66.800 ;
        RECT 76.400 66.800 78.200 67.600 ;
        RECT 79.600 66.800 81.800 67.600 ;
        RECT 82.800 66.800 85.000 67.600 ;
        RECT 86.000 66.800 88.400 67.600 ;
        RECT 90.800 67.400 91.400 70.400 ;
        RECT 92.600 69.600 93.200 71.800 ;
        RECT 94.000 71.800 95.400 72.400 ;
        RECT 96.000 71.800 97.000 72.400 ;
        RECT 100.400 71.800 101.200 79.800 ;
        RECT 102.000 72.400 102.800 79.800 ;
        RECT 105.200 72.400 106.000 79.800 ;
        RECT 102.000 71.800 106.000 72.400 ;
        RECT 94.000 71.600 94.800 71.800 ;
        RECT 89.200 66.800 91.400 67.400 ;
        RECT 76.400 62.200 77.200 66.800 ;
        RECT 79.600 62.200 80.400 66.800 ;
        RECT 82.800 62.200 83.600 66.800 ;
        RECT 86.000 62.200 86.800 66.800 ;
        RECT 89.200 62.200 90.000 66.800 ;
        RECT 92.400 62.200 93.200 69.600 ;
        RECT 96.000 68.400 96.600 71.800 ;
        RECT 100.600 70.400 101.200 71.800 ;
        RECT 106.800 71.400 107.600 79.800 ;
        RECT 111.200 76.400 112.000 79.800 ;
        RECT 110.000 75.800 112.000 76.400 ;
        RECT 115.600 75.800 116.400 79.800 ;
        RECT 119.800 75.800 121.000 79.800 ;
        RECT 110.000 75.000 110.800 75.800 ;
        RECT 115.600 75.200 116.200 75.800 ;
        RECT 113.400 74.600 117.000 75.200 ;
        RECT 119.600 75.000 120.400 75.800 ;
        RECT 113.400 74.400 114.200 74.600 ;
        RECT 116.200 74.400 117.000 74.600 ;
        RECT 124.400 74.300 125.200 79.800 ;
        RECT 126.000 74.300 126.800 74.400 ;
        RECT 110.000 73.000 110.800 73.200 ;
        RECT 114.600 73.000 115.400 73.200 ;
        RECT 110.000 72.400 115.400 73.000 ;
        RECT 116.000 73.000 118.200 73.600 ;
        RECT 116.000 71.800 116.600 73.000 ;
        RECT 117.400 72.800 118.200 73.000 ;
        RECT 119.800 73.200 121.200 74.000 ;
        RECT 124.400 73.700 126.800 74.300 ;
        RECT 119.800 72.200 120.400 73.200 ;
        RECT 111.800 71.400 116.600 71.800 ;
        RECT 106.800 71.200 116.600 71.400 ;
        RECT 118.000 71.600 120.400 72.200 ;
        RECT 106.800 71.000 112.600 71.200 ;
        RECT 106.800 70.800 112.400 71.000 ;
        RECT 104.400 70.400 105.200 70.800 ;
        RECT 97.200 68.800 98.000 70.400 ;
        RECT 100.400 69.800 102.800 70.400 ;
        RECT 104.400 69.800 106.000 70.400 ;
        RECT 113.200 70.200 114.000 70.400 ;
        RECT 100.400 69.600 101.200 69.800 ;
        RECT 102.200 68.400 102.800 69.800 ;
        RECT 105.200 69.600 106.000 69.800 ;
        RECT 109.000 69.600 114.000 70.200 ;
        RECT 109.000 69.400 109.800 69.600 ;
        RECT 111.600 69.400 112.400 69.600 ;
        RECT 94.000 67.600 96.600 68.400 ;
        RECT 98.800 68.200 99.600 68.400 ;
        RECT 98.000 67.600 99.600 68.200 ;
        RECT 102.000 67.600 102.800 68.400 ;
        RECT 103.600 68.300 104.400 69.200 ;
        RECT 110.600 68.400 111.400 68.600 ;
        RECT 118.000 68.400 118.600 71.600 ;
        RECT 124.400 71.200 125.200 73.700 ;
        RECT 126.000 73.600 126.800 73.700 ;
        RECT 121.000 70.600 125.200 71.200 ;
        RECT 121.000 70.400 121.800 70.600 ;
        RECT 122.600 69.800 123.400 70.000 ;
        RECT 119.600 69.200 123.400 69.800 ;
        RECT 119.600 69.000 120.400 69.200 ;
        RECT 105.200 68.300 106.000 68.400 ;
        RECT 103.600 67.700 106.000 68.300 ;
        RECT 103.600 67.600 104.400 67.700 ;
        RECT 105.200 67.600 106.000 67.700 ;
        RECT 107.600 67.800 118.600 68.400 ;
        RECT 107.600 67.600 109.200 67.800 ;
        RECT 94.200 66.200 94.800 67.600 ;
        RECT 98.000 67.200 98.800 67.600 ;
        RECT 95.800 66.200 99.400 66.600 ;
        RECT 94.000 62.200 94.800 66.200 ;
        RECT 95.600 66.000 99.600 66.200 ;
        RECT 95.600 62.200 96.400 66.000 ;
        RECT 98.800 62.200 99.600 66.000 ;
        RECT 100.400 65.600 101.200 66.400 ;
        RECT 102.200 66.200 102.800 67.600 ;
        RECT 100.600 64.800 101.400 65.600 ;
        RECT 102.000 62.200 102.800 66.200 ;
        RECT 106.800 62.200 107.600 67.000 ;
        RECT 111.800 65.600 112.400 67.800 ;
        RECT 117.400 67.600 118.200 67.800 ;
        RECT 124.400 67.200 125.200 70.600 ;
        RECT 121.400 66.600 125.200 67.200 ;
        RECT 121.400 66.400 122.200 66.600 ;
        RECT 110.000 64.200 110.800 65.000 ;
        RECT 111.600 64.800 112.400 65.600 ;
        RECT 113.400 65.400 114.200 65.600 ;
        RECT 113.400 64.800 116.200 65.400 ;
        RECT 115.600 64.200 116.200 64.800 ;
        RECT 119.600 64.200 120.400 65.000 ;
        RECT 110.000 63.600 112.000 64.200 ;
        RECT 111.200 62.200 112.000 63.600 ;
        RECT 115.600 62.200 116.400 64.200 ;
        RECT 119.600 63.600 121.000 64.200 ;
        RECT 119.800 62.200 121.000 63.600 ;
        RECT 124.400 62.200 125.200 66.600 ;
        RECT 127.600 68.300 128.400 79.800 ;
        RECT 131.800 72.400 132.600 79.800 ;
        RECT 142.000 75.800 142.800 79.800 ;
        RECT 133.200 73.600 134.000 74.400 ;
        RECT 133.400 72.400 134.000 73.600 ;
        RECT 131.800 71.800 132.800 72.400 ;
        RECT 133.400 71.800 134.800 72.400 ;
        RECT 130.800 68.800 131.600 70.400 ;
        RECT 132.200 70.300 132.800 71.800 ;
        RECT 134.000 71.600 134.800 71.800 ;
        RECT 142.200 71.600 142.800 75.800 ;
        RECT 145.200 71.800 146.000 79.800 ;
        RECT 142.200 71.000 144.600 71.600 ;
        RECT 138.800 70.300 139.600 70.400 ;
        RECT 132.200 69.700 139.600 70.300 ;
        RECT 132.200 68.400 132.800 69.700 ;
        RECT 138.800 69.600 139.600 69.700 ;
        RECT 142.000 69.600 142.800 70.400 ;
        RECT 129.200 68.300 130.000 68.400 ;
        RECT 127.600 68.200 130.000 68.300 ;
        RECT 127.600 67.700 130.800 68.200 ;
        RECT 126.000 64.800 126.800 66.400 ;
        RECT 127.600 62.200 128.400 67.700 ;
        RECT 129.200 67.600 130.800 67.700 ;
        RECT 132.200 67.600 134.800 68.400 ;
        RECT 140.400 67.600 141.200 69.200 ;
        RECT 142.200 68.800 142.800 69.600 ;
        RECT 142.200 68.200 143.200 68.800 ;
        RECT 142.400 68.000 143.200 68.200 ;
        RECT 144.000 67.600 144.600 71.000 ;
        RECT 145.400 70.400 146.000 71.800 ;
        RECT 145.200 69.600 146.000 70.400 ;
        RECT 130.000 67.200 130.800 67.600 ;
        RECT 129.400 66.200 133.000 66.600 ;
        RECT 134.000 66.200 134.600 67.600 ;
        RECT 144.000 67.400 144.800 67.600 ;
        RECT 141.800 67.000 144.800 67.400 ;
        RECT 140.600 66.800 144.800 67.000 ;
        RECT 140.600 66.400 142.400 66.800 ;
        RECT 140.600 66.200 141.200 66.400 ;
        RECT 145.400 66.200 146.000 69.600 ;
        RECT 129.200 66.000 133.200 66.200 ;
        RECT 129.200 62.200 130.000 66.000 ;
        RECT 132.400 62.200 133.200 66.000 ;
        RECT 134.000 62.200 134.800 66.200 ;
        RECT 140.400 62.200 141.200 66.200 ;
        RECT 144.600 65.200 146.000 66.200 ;
        RECT 144.600 62.200 145.400 65.200 ;
        RECT 146.800 62.200 147.600 79.800 ;
        RECT 150.000 68.300 150.800 68.400 ;
        RECT 148.500 67.700 150.800 68.300 ;
        RECT 148.500 66.400 149.100 67.700 ;
        RECT 150.000 66.800 150.800 67.700 ;
        RECT 148.400 64.800 149.200 66.400 ;
        RECT 151.600 66.200 152.400 79.800 ;
        RECT 153.200 71.600 154.000 73.200 ;
        RECT 154.800 71.200 155.600 79.800 ;
        RECT 159.000 75.800 160.200 79.800 ;
        RECT 163.600 75.800 164.400 79.800 ;
        RECT 168.000 76.400 168.800 79.800 ;
        RECT 168.000 75.800 170.000 76.400 ;
        RECT 159.600 75.000 160.400 75.800 ;
        RECT 163.800 75.200 164.400 75.800 ;
        RECT 163.000 74.600 166.600 75.200 ;
        RECT 169.200 75.000 170.000 75.800 ;
        RECT 163.000 74.400 163.800 74.600 ;
        RECT 165.800 74.400 166.600 74.600 ;
        RECT 158.800 73.200 160.200 74.000 ;
        RECT 159.600 72.200 160.200 73.200 ;
        RECT 161.800 73.000 164.000 73.600 ;
        RECT 161.800 72.800 162.600 73.000 ;
        RECT 159.600 71.600 162.000 72.200 ;
        RECT 154.800 70.600 159.000 71.200 ;
        RECT 154.800 67.200 155.600 70.600 ;
        RECT 158.200 70.400 159.000 70.600 ;
        RECT 156.600 69.800 157.400 70.000 ;
        RECT 156.600 69.200 160.400 69.800 ;
        RECT 159.600 69.000 160.400 69.200 ;
        RECT 161.400 68.400 162.000 71.600 ;
        RECT 163.400 71.800 164.000 73.000 ;
        RECT 164.600 73.000 165.400 73.200 ;
        RECT 169.200 73.000 170.000 73.200 ;
        RECT 164.600 72.400 170.000 73.000 ;
        RECT 163.400 71.400 168.200 71.800 ;
        RECT 172.400 71.400 173.200 79.800 ;
        RECT 163.400 71.200 173.200 71.400 ;
        RECT 167.400 71.000 173.200 71.200 ;
        RECT 167.600 70.800 173.200 71.000 ;
        RECT 174.000 71.400 174.800 79.800 ;
        RECT 178.400 76.400 179.200 79.800 ;
        RECT 177.200 75.800 179.200 76.400 ;
        RECT 182.800 75.800 183.600 79.800 ;
        RECT 187.000 75.800 188.200 79.800 ;
        RECT 177.200 75.000 178.000 75.800 ;
        RECT 182.800 75.200 183.400 75.800 ;
        RECT 180.600 74.600 184.200 75.200 ;
        RECT 186.800 75.000 187.600 75.800 ;
        RECT 180.600 74.400 181.400 74.600 ;
        RECT 183.400 74.400 184.200 74.600 ;
        RECT 177.200 73.000 178.000 73.200 ;
        RECT 181.800 73.000 182.600 73.200 ;
        RECT 177.200 72.400 182.600 73.000 ;
        RECT 183.200 73.000 185.400 73.600 ;
        RECT 183.200 71.800 183.800 73.000 ;
        RECT 184.600 72.800 185.400 73.000 ;
        RECT 187.000 73.200 188.400 74.000 ;
        RECT 187.000 72.200 187.600 73.200 ;
        RECT 179.000 71.400 183.800 71.800 ;
        RECT 174.000 71.200 183.800 71.400 ;
        RECT 185.200 71.600 187.600 72.200 ;
        RECT 174.000 71.000 179.800 71.200 ;
        RECT 174.000 70.800 179.600 71.000 ;
        RECT 166.000 70.200 166.800 70.400 ;
        RECT 180.400 70.200 181.200 70.400 ;
        RECT 166.000 69.600 171.000 70.200 ;
        RECT 170.200 69.400 171.000 69.600 ;
        RECT 176.200 69.600 181.200 70.200 ;
        RECT 176.200 69.400 177.000 69.600 ;
        RECT 178.800 69.400 179.600 69.600 ;
        RECT 168.600 68.400 169.400 68.600 ;
        RECT 177.800 68.400 178.600 68.600 ;
        RECT 185.200 68.400 185.800 71.600 ;
        RECT 191.600 71.200 192.400 79.800 ;
        RECT 188.200 70.600 192.400 71.200 ;
        RECT 188.200 70.400 189.000 70.600 ;
        RECT 189.800 69.800 190.600 70.000 ;
        RECT 186.800 69.200 190.600 69.800 ;
        RECT 186.800 69.000 187.600 69.200 ;
        RECT 161.400 67.800 172.400 68.400 ;
        RECT 161.800 67.600 162.600 67.800 ;
        RECT 154.800 66.600 158.600 67.200 ;
        RECT 151.600 65.600 153.400 66.200 ;
        RECT 152.600 64.400 153.400 65.600 ;
        RECT 152.600 63.600 154.000 64.400 ;
        RECT 152.600 62.200 153.400 63.600 ;
        RECT 154.800 62.200 155.600 66.600 ;
        RECT 157.800 66.400 158.600 66.600 ;
        RECT 167.600 66.400 168.200 67.800 ;
        RECT 170.800 67.600 172.400 67.800 ;
        RECT 174.800 67.800 185.800 68.400 ;
        RECT 174.800 67.600 176.400 67.800 ;
        RECT 165.800 65.400 166.600 65.600 ;
        RECT 159.600 64.200 160.400 65.000 ;
        RECT 163.800 64.800 166.600 65.400 ;
        RECT 167.600 64.800 168.400 66.400 ;
        RECT 163.800 64.200 164.400 64.800 ;
        RECT 169.200 64.200 170.000 65.000 ;
        RECT 159.000 63.600 160.400 64.200 ;
        RECT 159.000 62.200 160.200 63.600 ;
        RECT 163.600 62.200 164.400 64.200 ;
        RECT 168.000 63.600 170.000 64.200 ;
        RECT 168.000 62.200 168.800 63.600 ;
        RECT 172.400 62.200 173.200 67.000 ;
        RECT 174.000 62.200 174.800 67.000 ;
        RECT 179.000 65.600 179.600 67.800 ;
        RECT 184.600 67.600 185.400 67.800 ;
        RECT 191.600 67.200 192.400 70.600 ;
        RECT 188.600 66.600 192.400 67.200 ;
        RECT 188.600 66.400 189.400 66.600 ;
        RECT 177.200 64.200 178.000 65.000 ;
        RECT 178.800 64.800 179.600 65.600 ;
        RECT 180.600 65.400 181.400 65.600 ;
        RECT 180.600 64.800 183.400 65.400 ;
        RECT 182.800 64.200 183.400 64.800 ;
        RECT 186.800 64.200 187.600 65.000 ;
        RECT 177.200 63.600 179.200 64.200 ;
        RECT 178.400 62.200 179.200 63.600 ;
        RECT 182.800 62.200 183.600 64.200 ;
        RECT 186.800 63.600 188.200 64.200 ;
        RECT 187.000 62.200 188.200 63.600 ;
        RECT 191.600 62.200 192.400 66.600 ;
        RECT 4.400 55.200 5.200 59.800 ;
        RECT 3.000 54.600 5.200 55.200 ;
        RECT 6.000 55.400 6.800 59.800 ;
        RECT 10.200 58.400 11.400 59.800 ;
        RECT 10.200 57.800 11.600 58.400 ;
        RECT 14.800 57.800 15.600 59.800 ;
        RECT 19.200 58.400 20.000 59.800 ;
        RECT 19.200 57.800 21.200 58.400 ;
        RECT 10.800 57.000 11.600 57.800 ;
        RECT 15.000 57.200 15.600 57.800 ;
        RECT 15.000 56.600 17.800 57.200 ;
        RECT 17.000 56.400 17.800 56.600 ;
        RECT 18.800 56.400 19.600 57.200 ;
        RECT 20.400 57.000 21.200 57.800 ;
        RECT 9.000 55.400 9.800 55.600 ;
        RECT 6.000 54.800 9.800 55.400 ;
        RECT 3.000 51.600 3.600 54.600 ;
        RECT 4.400 52.300 5.200 53.200 ;
        RECT 6.000 52.300 6.800 54.800 ;
        RECT 13.000 54.200 13.800 54.400 ;
        RECT 17.200 54.200 18.000 54.400 ;
        RECT 18.800 54.200 19.400 56.400 ;
        RECT 23.600 55.000 24.400 59.800 ;
        RECT 25.200 55.800 26.000 59.800 ;
        RECT 29.400 58.400 30.200 59.800 ;
        RECT 29.400 57.600 30.800 58.400 ;
        RECT 29.400 56.800 30.200 57.600 ;
        RECT 29.400 55.800 30.800 56.800 ;
        RECT 25.400 55.600 26.000 55.800 ;
        RECT 25.400 55.200 27.200 55.600 ;
        RECT 25.400 55.000 29.600 55.200 ;
        RECT 26.600 54.600 29.600 55.000 ;
        RECT 28.800 54.400 29.600 54.600 ;
        RECT 22.000 54.200 23.600 54.400 ;
        RECT 12.600 53.600 23.600 54.200 ;
        RECT 10.800 52.800 11.600 53.000 ;
        RECT 4.400 51.700 6.800 52.300 ;
        RECT 7.800 52.200 11.600 52.800 ;
        RECT 7.800 52.000 8.600 52.200 ;
        RECT 4.400 51.600 5.200 51.700 ;
        RECT 2.400 50.800 3.600 51.600 ;
        RECT 3.000 50.200 3.600 50.800 ;
        RECT 6.000 51.400 6.800 51.700 ;
        RECT 9.400 51.400 10.200 51.600 ;
        RECT 6.000 50.800 10.200 51.400 ;
        RECT 3.000 49.600 5.200 50.200 ;
        RECT 4.400 42.200 5.200 49.600 ;
        RECT 6.000 42.200 6.800 50.800 ;
        RECT 12.600 50.400 13.200 53.600 ;
        RECT 19.800 53.400 20.600 53.600 ;
        RECT 26.800 53.200 28.000 54.000 ;
        RECT 18.800 52.400 19.600 52.600 ;
        RECT 21.400 52.400 22.200 52.600 ;
        RECT 27.000 52.400 27.600 53.200 ;
        RECT 17.200 51.800 22.200 52.400 ;
        RECT 17.200 51.600 18.000 51.800 ;
        RECT 26.800 51.600 27.600 52.400 ;
        RECT 18.800 51.000 24.400 51.200 ;
        RECT 28.800 51.000 29.400 54.400 ;
        RECT 30.200 52.400 30.800 55.800 ;
        RECT 33.200 55.200 34.000 59.800 ;
        RECT 36.400 55.200 37.200 59.800 ;
        RECT 39.600 55.200 40.400 59.800 ;
        RECT 42.800 55.200 43.600 59.800 ;
        RECT 30.000 51.600 30.800 52.400 ;
        RECT 18.600 50.800 24.400 51.000 ;
        RECT 10.800 49.800 13.200 50.400 ;
        RECT 14.600 50.600 24.400 50.800 ;
        RECT 14.600 50.200 19.400 50.600 ;
        RECT 10.800 48.800 11.400 49.800 ;
        RECT 10.000 48.000 11.400 48.800 ;
        RECT 13.000 49.000 13.800 49.200 ;
        RECT 14.600 49.000 15.200 50.200 ;
        RECT 13.000 48.400 15.200 49.000 ;
        RECT 15.800 49.000 21.200 49.600 ;
        RECT 15.800 48.800 16.600 49.000 ;
        RECT 20.400 48.800 21.200 49.000 ;
        RECT 14.200 47.400 15.000 47.600 ;
        RECT 17.000 47.400 17.800 47.600 ;
        RECT 10.800 46.200 11.600 47.000 ;
        RECT 14.200 46.800 17.800 47.400 ;
        RECT 15.000 46.200 15.600 46.800 ;
        RECT 20.400 46.200 21.200 47.000 ;
        RECT 10.200 42.200 11.400 46.200 ;
        RECT 14.800 42.200 15.600 46.200 ;
        RECT 19.200 45.600 21.200 46.200 ;
        RECT 19.200 42.200 20.000 45.600 ;
        RECT 23.600 42.200 24.400 50.600 ;
        RECT 27.000 50.400 29.400 51.000 ;
        RECT 27.000 46.200 27.600 50.400 ;
        RECT 30.200 50.200 30.800 51.600 ;
        RECT 31.600 54.400 34.000 55.200 ;
        RECT 35.000 54.400 37.200 55.200 ;
        RECT 38.200 54.400 40.400 55.200 ;
        RECT 41.800 54.400 43.600 55.200 ;
        RECT 50.800 55.000 51.600 59.800 ;
        RECT 55.200 58.400 56.000 59.800 ;
        RECT 54.000 57.800 56.000 58.400 ;
        RECT 59.600 57.800 60.400 59.800 ;
        RECT 63.800 58.400 65.000 59.800 ;
        RECT 63.600 57.800 65.000 58.400 ;
        RECT 54.000 57.000 54.800 57.800 ;
        RECT 59.600 57.200 60.200 57.800 ;
        RECT 55.600 56.400 56.400 57.200 ;
        RECT 57.400 56.600 60.200 57.200 ;
        RECT 63.600 57.000 64.400 57.800 ;
        RECT 57.400 56.400 58.200 56.600 ;
        RECT 31.600 51.600 32.400 54.400 ;
        RECT 35.000 53.800 35.800 54.400 ;
        RECT 38.200 53.800 39.000 54.400 ;
        RECT 41.800 53.800 42.600 54.400 ;
        RECT 33.200 53.000 35.800 53.800 ;
        RECT 36.600 53.000 39.000 53.800 ;
        RECT 40.000 53.000 42.600 53.800 ;
        RECT 51.600 54.200 53.200 54.400 ;
        RECT 55.800 54.200 56.400 56.400 ;
        RECT 65.400 55.400 66.200 55.600 ;
        RECT 68.400 55.400 69.200 59.800 ;
        RECT 72.600 56.400 73.400 59.800 ;
        RECT 76.400 57.800 77.200 59.800 ;
        RECT 65.400 54.800 69.200 55.400 ;
        RECT 71.600 56.300 73.400 56.400 ;
        RECT 74.800 56.300 75.600 57.200 ;
        RECT 71.600 55.700 75.600 56.300 ;
        RECT 61.400 54.200 62.200 54.400 ;
        RECT 51.600 53.600 62.600 54.200 ;
        RECT 54.600 53.400 55.400 53.600 ;
        RECT 35.000 51.600 35.800 53.000 ;
        RECT 38.200 51.600 39.000 53.000 ;
        RECT 41.800 51.600 42.600 53.000 ;
        RECT 53.000 52.400 53.800 52.600 ;
        RECT 53.000 51.800 58.000 52.400 ;
        RECT 57.200 51.600 58.000 51.800 ;
        RECT 31.600 50.800 34.000 51.600 ;
        RECT 35.000 50.800 37.200 51.600 ;
        RECT 38.200 50.800 40.400 51.600 ;
        RECT 41.800 50.800 43.600 51.600 ;
        RECT 26.800 42.200 27.600 46.200 ;
        RECT 30.000 42.200 30.800 50.200 ;
        RECT 33.200 42.200 34.000 50.800 ;
        RECT 36.400 42.200 37.200 50.800 ;
        RECT 39.600 42.200 40.400 50.800 ;
        RECT 42.800 42.200 43.600 50.800 ;
        RECT 50.800 51.000 56.400 51.200 ;
        RECT 50.800 50.800 56.600 51.000 ;
        RECT 50.800 50.600 60.600 50.800 ;
        RECT 50.800 42.200 51.600 50.600 ;
        RECT 55.800 50.200 60.600 50.600 ;
        RECT 54.000 49.000 59.400 49.600 ;
        RECT 54.000 48.800 54.800 49.000 ;
        RECT 58.600 48.800 59.400 49.000 ;
        RECT 60.000 49.000 60.600 50.200 ;
        RECT 62.000 50.400 62.600 53.600 ;
        RECT 63.600 52.800 64.400 53.000 ;
        RECT 63.600 52.200 67.400 52.800 ;
        RECT 66.600 52.000 67.400 52.200 ;
        RECT 65.000 51.400 65.800 51.600 ;
        RECT 68.400 51.400 69.200 54.800 ;
        RECT 70.000 53.600 70.800 55.200 ;
        RECT 65.000 50.800 69.200 51.400 ;
        RECT 62.000 49.800 64.400 50.400 ;
        RECT 61.400 49.000 62.200 49.200 ;
        RECT 60.000 48.400 62.200 49.000 ;
        RECT 63.800 48.800 64.400 49.800 ;
        RECT 63.800 48.000 65.200 48.800 ;
        RECT 57.400 47.400 58.200 47.600 ;
        RECT 60.200 47.400 61.000 47.600 ;
        RECT 54.000 46.200 54.800 47.000 ;
        RECT 57.400 46.800 61.000 47.400 ;
        RECT 59.600 46.200 60.200 46.800 ;
        RECT 63.600 46.200 64.400 47.000 ;
        RECT 54.000 45.600 56.000 46.200 ;
        RECT 55.200 42.200 56.000 45.600 ;
        RECT 59.600 42.200 60.400 46.200 ;
        RECT 63.800 42.200 65.000 46.200 ;
        RECT 68.400 42.200 69.200 50.800 ;
        RECT 71.600 42.200 72.400 55.700 ;
        RECT 74.800 55.600 75.600 55.700 ;
        RECT 76.600 54.400 77.200 57.800 ;
        RECT 79.800 56.400 80.600 57.200 ;
        RECT 79.600 55.600 80.400 56.400 ;
        RECT 81.200 55.800 82.000 59.800 ;
        RECT 88.600 56.400 89.400 59.800 ;
        RECT 76.400 53.600 77.200 54.400 ;
        RECT 73.200 52.300 74.000 52.400 ;
        RECT 76.600 52.300 77.200 53.600 ;
        RECT 73.200 51.700 77.200 52.300 ;
        RECT 73.200 51.600 74.000 51.700 ;
        RECT 73.200 48.800 74.000 50.400 ;
        RECT 76.600 50.200 77.200 51.700 ;
        RECT 78.000 52.300 78.800 52.400 ;
        RECT 79.600 52.300 80.400 52.400 ;
        RECT 78.000 52.200 80.400 52.300 ;
        RECT 81.400 52.200 82.000 55.800 ;
        RECT 87.600 55.600 90.000 56.400 ;
        RECT 82.800 52.800 83.600 54.400 ;
        RECT 86.000 53.600 86.800 55.200 ;
        RECT 84.400 52.200 85.200 52.400 ;
        RECT 78.000 51.700 82.000 52.200 ;
        RECT 78.000 50.800 78.800 51.700 ;
        RECT 79.600 51.600 82.000 51.700 ;
        RECT 83.600 51.600 85.200 52.200 ;
        RECT 79.800 50.200 80.400 51.600 ;
        RECT 83.600 51.200 84.400 51.600 ;
        RECT 76.400 49.400 78.200 50.200 ;
        RECT 77.400 42.200 78.200 49.400 ;
        RECT 79.600 42.200 80.400 50.200 ;
        RECT 81.200 49.600 85.200 50.200 ;
        RECT 81.200 42.200 82.000 49.600 ;
        RECT 84.400 42.200 85.200 49.600 ;
        RECT 87.600 42.200 88.400 55.600 ;
        RECT 92.400 55.200 93.200 59.800 ;
        RECT 95.600 55.200 96.400 59.800 ;
        RECT 98.800 55.200 99.600 59.800 ;
        RECT 102.000 55.200 102.800 59.800 ;
        RECT 105.800 58.400 106.600 59.800 ;
        RECT 105.200 57.600 106.600 58.400 ;
        RECT 111.600 57.800 112.400 59.800 ;
        RECT 119.600 57.800 120.400 59.800 ;
        RECT 122.800 58.400 123.600 59.800 ;
        RECT 105.800 56.400 106.600 57.600 ;
        RECT 105.800 55.800 107.600 56.400 ;
        RECT 92.400 54.400 94.200 55.200 ;
        RECT 95.600 54.400 97.800 55.200 ;
        RECT 98.800 54.400 101.000 55.200 ;
        RECT 102.000 54.400 104.400 55.200 ;
        RECT 93.400 53.800 94.200 54.400 ;
        RECT 97.000 53.800 97.800 54.400 ;
        RECT 100.200 53.800 101.000 54.400 ;
        RECT 93.400 53.000 96.000 53.800 ;
        RECT 97.000 53.000 99.400 53.800 ;
        RECT 100.200 53.000 102.800 53.800 ;
        RECT 93.400 51.600 94.200 53.000 ;
        RECT 97.000 51.600 97.800 53.000 ;
        RECT 100.200 51.600 101.000 53.000 ;
        RECT 103.600 51.600 104.400 54.400 ;
        RECT 92.400 50.800 94.200 51.600 ;
        RECT 95.600 50.800 97.800 51.600 ;
        RECT 98.800 50.800 101.000 51.600 ;
        RECT 102.000 50.800 104.400 51.600 ;
        RECT 89.200 48.800 90.000 50.400 ;
        RECT 92.400 42.200 93.200 50.800 ;
        RECT 95.600 42.200 96.400 50.800 ;
        RECT 98.800 42.200 99.600 50.800 ;
        RECT 102.000 42.200 102.800 50.800 ;
        RECT 105.200 48.800 106.000 50.400 ;
        RECT 106.800 42.200 107.600 55.800 ;
        RECT 110.000 55.600 110.800 57.200 ;
        RECT 108.400 54.300 109.200 55.200 ;
        RECT 111.800 54.400 112.400 57.800 ;
        RECT 119.200 57.600 120.400 57.800 ;
        RECT 122.600 57.600 123.600 58.400 ;
        RECT 119.200 57.000 123.200 57.600 ;
        RECT 111.600 54.300 112.400 54.400 ;
        RECT 116.400 54.300 117.200 54.400 ;
        RECT 108.400 53.700 117.200 54.300 ;
        RECT 108.400 53.600 109.200 53.700 ;
        RECT 111.600 53.600 112.400 53.700 ;
        RECT 116.400 53.600 117.200 53.700 ;
        RECT 111.800 50.200 112.400 53.600 ;
        RECT 113.200 52.300 114.000 52.400 ;
        RECT 116.400 52.300 117.200 52.400 ;
        RECT 113.200 51.700 117.200 52.300 ;
        RECT 113.200 50.800 114.000 51.700 ;
        RECT 116.400 51.600 117.200 51.700 ;
        RECT 119.200 50.400 119.800 57.000 ;
        RECT 122.800 55.600 125.200 56.400 ;
        RECT 127.600 56.000 128.400 59.800 ;
        RECT 130.800 56.000 131.600 59.800 ;
        RECT 127.600 55.800 131.600 56.000 ;
        RECT 132.400 55.800 133.200 59.800 ;
        RECT 139.400 58.400 140.200 59.800 ;
        RECT 138.800 57.600 140.200 58.400 ;
        RECT 139.400 56.800 140.200 57.600 ;
        RECT 138.800 55.800 140.200 56.800 ;
        RECT 143.600 55.800 144.400 59.800 ;
        RECT 145.800 58.400 146.600 59.800 ;
        RECT 145.200 57.600 146.600 58.400 ;
        RECT 145.800 56.400 146.600 57.600 ;
        RECT 145.800 55.800 147.600 56.400 ;
        RECT 150.000 55.800 150.800 59.800 ;
        RECT 154.200 56.800 155.000 59.800 ;
        RECT 154.200 55.800 155.600 56.800 ;
        RECT 127.800 55.400 131.400 55.800 ;
        RECT 128.400 54.400 129.200 54.800 ;
        RECT 132.400 54.400 133.000 55.800 ;
        RECT 122.000 54.300 123.600 54.400 ;
        RECT 127.600 54.300 129.200 54.400 ;
        RECT 122.000 53.800 129.200 54.300 ;
        RECT 122.000 53.700 128.400 53.800 ;
        RECT 122.000 53.600 123.600 53.700 ;
        RECT 127.600 53.600 128.400 53.700 ;
        RECT 130.600 53.600 133.200 54.400 ;
        RECT 120.400 51.600 122.000 52.400 ;
        RECT 129.200 51.600 130.000 53.200 ;
        RECT 111.600 49.400 113.400 50.200 ;
        RECT 116.400 49.800 119.800 50.400 ;
        RECT 130.600 50.200 131.200 53.600 ;
        RECT 138.800 52.400 139.400 55.800 ;
        RECT 143.600 55.600 144.200 55.800 ;
        RECT 142.400 55.200 144.200 55.600 ;
        RECT 140.000 55.000 144.200 55.200 ;
        RECT 140.000 54.600 143.000 55.000 ;
        RECT 140.000 54.400 140.800 54.600 ;
        RECT 138.800 51.600 139.600 52.400 ;
        RECT 132.400 50.200 133.200 50.400 ;
        RECT 116.400 49.600 117.200 49.800 ;
        RECT 112.600 42.200 113.400 49.400 ;
        RECT 116.600 49.000 117.200 49.600 ;
        RECT 130.200 49.600 131.200 50.200 ;
        RECT 131.800 49.600 133.200 50.200 ;
        RECT 138.800 50.200 139.400 51.600 ;
        RECT 140.200 51.000 140.800 54.400 ;
        RECT 141.600 53.800 142.400 54.000 ;
        RECT 141.600 53.200 142.600 53.800 ;
        RECT 142.000 52.400 142.600 53.200 ;
        RECT 143.600 52.800 144.400 54.400 ;
        RECT 142.000 51.600 142.800 52.400 ;
        RECT 140.200 50.400 142.600 51.000 ;
        RECT 118.200 49.000 121.800 49.200 ;
        RECT 114.800 43.000 115.600 49.000 ;
        RECT 116.400 43.400 117.200 49.000 ;
        RECT 118.000 48.600 121.800 49.000 ;
        RECT 115.000 42.800 115.600 43.000 ;
        RECT 118.000 43.000 118.800 48.600 ;
        RECT 121.200 48.200 121.800 48.600 ;
        RECT 123.000 48.800 126.600 49.400 ;
        RECT 123.000 48.200 123.600 48.800 ;
        RECT 118.000 42.800 118.600 43.000 ;
        RECT 115.000 42.200 118.600 42.800 ;
        RECT 119.600 42.800 120.400 48.000 ;
        RECT 121.200 43.400 122.000 48.200 ;
        RECT 122.800 42.800 123.600 48.200 ;
        RECT 119.600 42.200 123.600 42.800 ;
        RECT 126.000 48.200 126.600 48.800 ;
        RECT 126.000 42.200 126.800 48.200 ;
        RECT 130.200 44.400 131.000 49.600 ;
        RECT 131.800 48.400 132.400 49.600 ;
        RECT 131.600 47.600 132.400 48.400 ;
        RECT 129.200 43.600 131.000 44.400 ;
        RECT 130.200 42.200 131.000 43.600 ;
        RECT 138.800 42.200 139.600 50.200 ;
        RECT 142.000 46.200 142.600 50.400 ;
        RECT 145.200 48.800 146.000 50.400 ;
        RECT 142.000 42.200 142.800 46.200 ;
        RECT 146.800 42.200 147.600 55.800 ;
        RECT 150.200 55.600 150.800 55.800 ;
        RECT 150.200 55.200 152.000 55.600 ;
        RECT 148.400 53.600 149.200 55.200 ;
        RECT 150.200 55.000 154.400 55.200 ;
        RECT 151.400 54.600 154.400 55.000 ;
        RECT 153.600 54.400 154.400 54.600 ;
        RECT 150.000 52.800 150.800 54.400 ;
        RECT 152.000 53.800 152.800 54.000 ;
        RECT 151.800 53.200 152.800 53.800 ;
        RECT 151.800 52.400 152.400 53.200 ;
        RECT 151.600 51.600 152.400 52.400 ;
        RECT 153.600 51.000 154.200 54.400 ;
        RECT 155.000 52.400 155.600 55.800 ;
        RECT 158.000 56.300 158.800 56.400 ;
        RECT 160.000 56.300 160.800 59.800 ;
        RECT 158.000 55.700 160.800 56.300 ;
        RECT 158.000 55.600 158.800 55.700 ;
        RECT 160.000 54.200 160.800 55.700 ;
        RECT 164.000 58.400 164.800 59.800 ;
        RECT 164.000 57.600 165.200 58.400 ;
        RECT 170.800 57.800 171.600 59.800 ;
        RECT 174.600 58.400 175.400 59.800 ;
        RECT 164.000 54.200 164.800 57.600 ;
        RECT 169.200 55.600 170.000 57.200 ;
        RECT 171.000 54.400 171.600 57.800 ;
        RECT 174.000 57.600 175.400 58.400 ;
        RECT 174.600 56.800 175.400 57.600 ;
        RECT 160.000 53.800 161.800 54.200 ;
        RECT 160.200 53.600 161.800 53.800 ;
        RECT 154.800 51.600 155.600 52.400 ;
        RECT 158.000 51.600 159.600 52.400 ;
        RECT 151.800 50.400 154.200 51.000 ;
        RECT 155.000 50.400 155.600 51.600 ;
        RECT 151.800 46.200 152.400 50.400 ;
        RECT 151.600 42.200 152.400 46.200 ;
        RECT 154.800 50.300 155.600 50.400 ;
        RECT 156.400 50.300 157.200 51.200 ;
        RECT 154.800 49.700 157.200 50.300 ;
        RECT 154.800 42.200 155.600 49.700 ;
        RECT 156.400 49.600 157.200 49.700 ;
        RECT 161.200 50.400 161.800 53.600 ;
        RECT 163.000 53.800 164.800 54.200 ;
        RECT 163.000 53.600 164.600 53.800 ;
        RECT 170.800 53.600 171.600 54.400 ;
        RECT 163.000 50.400 163.600 53.600 ;
        RECT 165.200 51.600 166.800 52.400 ;
        RECT 169.200 52.300 170.000 52.400 ;
        RECT 171.000 52.300 171.600 53.600 ;
        RECT 174.000 55.800 175.400 56.800 ;
        RECT 178.800 55.800 179.600 59.800 ;
        RECT 181.000 56.400 181.800 59.800 ;
        RECT 174.000 52.400 174.600 55.800 ;
        RECT 178.800 55.600 179.400 55.800 ;
        RECT 180.400 55.600 182.800 56.400 ;
        RECT 177.600 55.200 179.400 55.600 ;
        RECT 175.200 55.000 179.400 55.200 ;
        RECT 175.200 54.600 178.200 55.000 ;
        RECT 175.200 54.400 176.000 54.600 ;
        RECT 169.200 51.700 171.600 52.300 ;
        RECT 169.200 51.600 170.000 51.700 ;
        RECT 161.200 49.600 162.000 50.400 ;
        RECT 162.800 49.600 163.600 50.400 ;
        RECT 167.600 49.600 168.400 51.200 ;
        RECT 171.000 50.200 171.600 51.700 ;
        RECT 172.400 50.800 173.200 52.400 ;
        RECT 174.000 51.600 174.800 52.400 ;
        RECT 174.000 50.200 174.600 51.600 ;
        RECT 175.400 51.000 176.000 54.400 ;
        RECT 178.800 54.300 179.600 54.400 ;
        RECT 180.400 54.300 181.200 54.400 ;
        RECT 176.800 53.800 177.600 54.000 ;
        RECT 176.800 53.200 177.800 53.800 ;
        RECT 177.200 52.400 177.800 53.200 ;
        RECT 178.800 53.700 181.200 54.300 ;
        RECT 178.800 52.800 179.600 53.700 ;
        RECT 180.400 53.600 181.200 53.700 ;
        RECT 177.200 51.600 178.000 52.400 ;
        RECT 175.400 50.400 177.800 51.000 ;
        RECT 158.000 48.300 158.800 48.400 ;
        RECT 159.600 48.300 160.400 49.200 ;
        RECT 158.000 47.700 160.400 48.300 ;
        RECT 158.000 47.600 158.800 47.700 ;
        RECT 159.600 47.600 160.400 47.700 ;
        RECT 161.200 47.000 161.800 49.600 ;
        RECT 158.200 46.400 161.800 47.000 ;
        RECT 158.200 46.200 158.800 46.400 ;
        RECT 158.000 42.200 158.800 46.200 ;
        RECT 161.200 46.200 161.800 46.400 ;
        RECT 163.000 47.000 163.600 49.600 ;
        RECT 170.800 49.400 172.600 50.200 ;
        RECT 164.400 47.600 165.200 49.200 ;
        RECT 163.000 46.400 166.600 47.000 ;
        RECT 163.000 46.200 163.600 46.400 ;
        RECT 161.200 42.200 162.000 46.200 ;
        RECT 162.800 42.200 163.600 46.200 ;
        RECT 166.000 46.200 166.600 46.400 ;
        RECT 166.000 42.200 166.800 46.200 ;
        RECT 171.800 42.200 172.600 49.400 ;
        RECT 174.000 42.200 174.800 50.200 ;
        RECT 177.200 46.200 177.800 50.400 ;
        RECT 178.800 50.300 179.600 50.400 ;
        RECT 180.400 50.300 181.200 50.400 ;
        RECT 178.800 49.700 181.200 50.300 ;
        RECT 178.800 49.600 179.600 49.700 ;
        RECT 180.400 48.800 181.200 49.700 ;
        RECT 177.200 42.200 178.000 46.200 ;
        RECT 182.000 42.200 182.800 55.600 ;
        RECT 185.200 55.200 186.000 59.800 ;
        RECT 190.000 55.200 190.800 59.800 ;
        RECT 183.600 53.600 184.400 55.200 ;
        RECT 185.200 54.600 187.400 55.200 ;
        RECT 190.000 54.600 192.200 55.200 ;
        RECT 183.700 52.300 184.300 53.600 ;
        RECT 185.200 52.300 186.000 53.200 ;
        RECT 183.700 51.700 186.000 52.300 ;
        RECT 185.200 51.600 186.000 51.700 ;
        RECT 186.800 51.600 187.400 54.600 ;
        RECT 190.000 51.600 190.800 53.200 ;
        RECT 191.600 51.600 192.200 54.600 ;
        RECT 186.800 50.800 188.000 51.600 ;
        RECT 191.600 50.800 192.800 51.600 ;
        RECT 186.800 50.200 187.400 50.800 ;
        RECT 191.600 50.200 192.200 50.800 ;
        RECT 185.200 49.600 187.400 50.200 ;
        RECT 190.000 49.600 192.200 50.200 ;
        RECT 185.200 42.200 186.000 49.600 ;
        RECT 190.000 42.200 190.800 49.600 ;
        RECT 1.200 31.200 2.000 39.800 ;
        RECT 5.400 35.800 6.600 39.800 ;
        RECT 10.000 35.800 10.800 39.800 ;
        RECT 14.400 36.400 15.200 39.800 ;
        RECT 14.400 35.800 16.400 36.400 ;
        RECT 6.000 35.000 6.800 35.800 ;
        RECT 10.200 35.200 10.800 35.800 ;
        RECT 9.400 34.600 13.000 35.200 ;
        RECT 15.600 35.000 16.400 35.800 ;
        RECT 9.400 34.400 10.200 34.600 ;
        RECT 12.200 34.400 13.000 34.600 ;
        RECT 5.200 33.200 6.600 34.000 ;
        RECT 6.000 32.200 6.600 33.200 ;
        RECT 8.200 33.000 10.400 33.600 ;
        RECT 8.200 32.800 9.000 33.000 ;
        RECT 6.000 31.600 8.400 32.200 ;
        RECT 1.200 30.600 5.400 31.200 ;
        RECT 1.200 27.200 2.000 30.600 ;
        RECT 4.600 30.400 5.400 30.600 ;
        RECT 3.000 29.800 3.800 30.000 ;
        RECT 3.000 29.200 6.800 29.800 ;
        RECT 6.000 29.000 6.800 29.200 ;
        RECT 7.800 28.400 8.400 31.600 ;
        RECT 9.800 31.800 10.400 33.000 ;
        RECT 11.000 33.000 11.800 33.200 ;
        RECT 15.600 33.000 16.400 33.200 ;
        RECT 11.000 32.400 16.400 33.000 ;
        RECT 9.800 31.400 14.600 31.800 ;
        RECT 18.800 31.400 19.600 39.800 ;
        RECT 21.200 33.600 22.000 34.400 ;
        RECT 21.200 32.400 21.800 33.600 ;
        RECT 22.600 32.400 23.400 39.800 ;
        RECT 29.400 32.600 30.200 39.800 ;
        RECT 20.400 31.800 21.800 32.400 ;
        RECT 22.400 31.800 23.400 32.400 ;
        RECT 28.400 31.800 30.200 32.600 ;
        RECT 32.400 33.600 33.200 34.400 ;
        RECT 32.400 32.400 33.000 33.600 ;
        RECT 33.800 32.400 34.600 39.800 ;
        RECT 31.600 31.800 33.000 32.400 ;
        RECT 33.600 31.800 34.600 32.400 ;
        RECT 20.400 31.600 21.200 31.800 ;
        RECT 9.800 31.200 19.600 31.400 ;
        RECT 13.800 31.000 19.600 31.200 ;
        RECT 14.000 30.800 19.600 31.000 ;
        RECT 12.400 30.200 13.200 30.400 ;
        RECT 12.400 29.600 17.400 30.200 ;
        RECT 14.000 29.400 14.800 29.600 ;
        RECT 16.600 29.400 17.400 29.600 ;
        RECT 15.000 28.400 15.800 28.600 ;
        RECT 22.400 28.400 23.000 31.800 ;
        RECT 23.600 28.800 24.400 30.400 ;
        RECT 25.200 30.300 26.000 30.400 ;
        RECT 28.600 30.300 29.200 31.800 ;
        RECT 31.600 31.600 32.400 31.800 ;
        RECT 25.200 29.700 29.200 30.300 ;
        RECT 25.200 29.600 26.000 29.700 ;
        RECT 28.600 28.400 29.200 29.700 ;
        RECT 30.000 30.300 30.800 31.200 ;
        RECT 33.600 30.300 34.200 31.800 ;
        RECT 30.000 29.700 34.200 30.300 ;
        RECT 30.000 29.600 30.800 29.700 ;
        RECT 33.600 28.400 34.200 29.700 ;
        RECT 7.800 27.800 18.800 28.400 ;
        RECT 8.200 27.600 9.000 27.800 ;
        RECT 1.200 26.600 5.000 27.200 ;
        RECT 1.200 22.200 2.000 26.600 ;
        RECT 4.200 26.400 5.000 26.600 ;
        RECT 14.000 25.600 14.600 27.800 ;
        RECT 17.200 27.600 18.800 27.800 ;
        RECT 20.400 27.600 23.000 28.400 ;
        RECT 25.200 28.200 26.000 28.400 ;
        RECT 24.400 27.600 26.000 28.200 ;
        RECT 28.400 27.600 29.200 28.400 ;
        RECT 31.600 27.600 34.200 28.400 ;
        RECT 36.400 28.300 37.200 28.400 ;
        RECT 38.000 28.300 38.800 28.400 ;
        RECT 36.400 28.200 38.800 28.300 ;
        RECT 35.600 27.700 38.800 28.200 ;
        RECT 35.600 27.600 37.200 27.700 ;
        RECT 12.200 25.400 13.000 25.600 ;
        RECT 6.000 24.200 6.800 25.000 ;
        RECT 10.200 24.800 13.000 25.400 ;
        RECT 14.000 24.800 14.800 25.600 ;
        RECT 10.200 24.200 10.800 24.800 ;
        RECT 15.600 24.200 16.400 25.000 ;
        RECT 5.400 23.600 6.800 24.200 ;
        RECT 5.400 22.200 6.600 23.600 ;
        RECT 10.000 22.200 10.800 24.200 ;
        RECT 14.400 23.600 16.400 24.200 ;
        RECT 14.400 22.200 15.200 23.600 ;
        RECT 18.800 22.200 19.600 27.000 ;
        RECT 20.600 26.200 21.200 27.600 ;
        RECT 24.400 27.200 25.200 27.600 ;
        RECT 22.200 26.200 25.800 26.600 ;
        RECT 20.400 22.200 21.200 26.200 ;
        RECT 22.000 26.000 26.000 26.200 ;
        RECT 22.000 22.200 22.800 26.000 ;
        RECT 25.200 22.200 26.000 26.000 ;
        RECT 26.800 24.800 27.600 26.400 ;
        RECT 28.600 24.200 29.200 27.600 ;
        RECT 31.800 26.200 32.400 27.600 ;
        RECT 35.600 27.200 36.400 27.600 ;
        RECT 38.000 26.800 38.800 27.700 ;
        RECT 39.600 28.300 40.400 39.800 ;
        RECT 43.600 33.600 44.400 34.400 ;
        RECT 43.600 32.400 44.200 33.600 ;
        RECT 45.000 32.400 45.800 39.800 ;
        RECT 51.800 32.600 52.600 39.800 ;
        RECT 42.800 31.800 44.200 32.400 ;
        RECT 44.800 31.800 45.800 32.400 ;
        RECT 50.800 31.800 52.600 32.600 ;
        RECT 42.800 31.600 43.600 31.800 ;
        RECT 44.800 28.400 45.400 31.800 ;
        RECT 46.000 28.800 46.800 30.400 ;
        RECT 51.000 28.400 51.600 31.800 ;
        RECT 58.800 31.600 59.600 33.200 ;
        RECT 52.400 30.300 53.200 31.200 ;
        RECT 60.400 30.300 61.200 39.800 ;
        RECT 65.200 35.800 66.000 39.800 ;
        RECT 65.400 31.600 66.000 35.800 ;
        RECT 68.400 31.800 69.200 39.800 ;
        RECT 70.000 35.800 70.800 39.800 ;
        RECT 70.200 35.600 70.800 35.800 ;
        RECT 73.200 35.800 74.000 39.800 ;
        RECT 73.200 35.600 73.800 35.800 ;
        RECT 70.200 35.000 73.800 35.600 ;
        RECT 70.200 32.400 70.800 35.000 ;
        RECT 71.600 32.800 72.400 34.400 ;
        RECT 65.400 31.000 67.800 31.600 ;
        RECT 52.400 29.700 61.200 30.300 ;
        RECT 52.400 29.600 53.200 29.700 ;
        RECT 41.200 28.300 42.000 28.400 ;
        RECT 39.600 27.700 42.000 28.300 ;
        RECT 33.400 26.200 37.000 26.600 ;
        RECT 39.600 26.200 40.400 27.700 ;
        RECT 41.200 27.600 42.000 27.700 ;
        RECT 42.800 27.600 45.400 28.400 ;
        RECT 47.600 28.300 48.400 28.400 ;
        RECT 50.800 28.300 51.600 28.400 ;
        RECT 58.800 28.300 59.600 28.400 ;
        RECT 47.600 28.200 49.900 28.300 ;
        RECT 46.800 27.700 49.900 28.200 ;
        RECT 46.800 27.600 48.400 27.700 ;
        RECT 43.000 26.200 43.600 27.600 ;
        RECT 46.800 27.200 47.600 27.600 ;
        RECT 44.600 26.200 48.200 26.600 ;
        RECT 49.300 26.400 49.900 27.700 ;
        RECT 50.800 27.700 59.600 28.300 ;
        RECT 50.800 27.600 51.600 27.700 ;
        RECT 58.800 27.600 59.600 27.700 ;
        RECT 28.400 22.200 29.200 24.200 ;
        RECT 31.600 22.200 32.400 26.200 ;
        RECT 33.200 26.000 37.200 26.200 ;
        RECT 33.200 22.200 34.000 26.000 ;
        RECT 36.400 22.200 37.200 26.000 ;
        RECT 39.600 25.600 41.400 26.200 ;
        RECT 40.600 22.200 41.400 25.600 ;
        RECT 42.800 22.200 43.600 26.200 ;
        RECT 44.400 26.000 48.400 26.200 ;
        RECT 44.400 22.200 45.200 26.000 ;
        RECT 47.600 22.200 48.400 26.000 ;
        RECT 49.200 24.800 50.000 26.400 ;
        RECT 51.000 24.200 51.600 27.600 ;
        RECT 60.400 26.200 61.200 29.700 ;
        RECT 65.200 29.600 66.000 30.400 ;
        RECT 62.000 28.300 62.800 28.400 ;
        RECT 63.600 28.300 64.400 29.200 ;
        RECT 62.000 27.700 64.400 28.300 ;
        RECT 65.400 28.800 66.000 29.600 ;
        RECT 65.400 28.200 66.400 28.800 ;
        RECT 65.600 28.000 66.400 28.200 ;
        RECT 62.000 26.800 62.800 27.700 ;
        RECT 63.600 27.600 64.400 27.700 ;
        RECT 67.200 27.600 67.800 31.000 ;
        RECT 68.600 30.400 69.200 31.800 ;
        RECT 70.000 31.600 70.800 32.400 ;
        RECT 68.400 29.600 69.200 30.400 ;
        RECT 67.200 27.400 68.000 27.600 ;
        RECT 65.000 27.000 68.000 27.400 ;
        RECT 63.800 26.800 68.000 27.000 ;
        RECT 63.800 26.400 65.600 26.800 ;
        RECT 63.800 26.200 64.400 26.400 ;
        RECT 68.600 26.200 69.200 29.600 ;
        RECT 70.200 28.400 70.800 31.600 ;
        RECT 74.800 32.300 75.600 32.400 ;
        RECT 76.400 32.300 77.200 39.800 ;
        RECT 74.800 31.800 77.200 32.300 ;
        RECT 79.600 35.800 80.400 39.800 ;
        RECT 74.800 31.700 77.100 31.800 ;
        RECT 74.800 30.800 75.600 31.700 ;
        RECT 76.400 30.400 77.000 31.700 ;
        RECT 79.600 31.600 80.200 35.800 ;
        RECT 82.800 32.400 83.600 39.800 ;
        RECT 86.000 32.400 86.800 39.800 ;
        RECT 82.800 31.800 86.800 32.400 ;
        RECT 87.600 31.800 88.400 39.800 ;
        RECT 91.800 32.400 92.600 39.800 ;
        RECT 93.200 33.600 94.000 34.400 ;
        RECT 93.400 32.400 94.000 33.600 ;
        RECT 96.400 33.600 97.200 34.400 ;
        RECT 96.400 32.400 97.000 33.600 ;
        RECT 97.800 32.400 98.600 39.800 ;
        RECT 91.800 31.800 92.800 32.400 ;
        RECT 93.400 32.300 94.800 32.400 ;
        RECT 95.600 32.300 97.000 32.400 ;
        RECT 93.400 31.800 97.000 32.300 ;
        RECT 97.600 31.800 98.600 32.400 ;
        RECT 102.000 32.400 102.800 39.800 ;
        RECT 105.200 32.400 106.000 39.800 ;
        RECT 102.000 31.800 106.000 32.400 ;
        RECT 106.800 31.800 107.600 39.800 ;
        RECT 77.800 31.000 80.200 31.600 ;
        RECT 72.400 29.600 74.000 30.400 ;
        RECT 76.400 29.600 77.200 30.400 ;
        RECT 70.200 28.200 71.800 28.400 ;
        RECT 70.200 27.800 72.000 28.200 ;
        RECT 50.800 22.200 51.600 24.200 ;
        RECT 59.400 25.600 61.200 26.200 ;
        RECT 59.400 22.200 60.200 25.600 ;
        RECT 63.600 22.200 64.400 26.200 ;
        RECT 67.800 25.200 69.200 26.200 ;
        RECT 67.800 22.200 68.600 25.200 ;
        RECT 71.200 22.200 72.000 27.800 ;
        RECT 76.400 26.200 77.000 29.600 ;
        RECT 77.800 27.600 78.400 31.000 ;
        RECT 83.600 30.400 84.400 30.800 ;
        RECT 87.600 30.400 88.200 31.800 ;
        RECT 79.600 29.600 80.400 30.400 ;
        RECT 82.800 29.800 84.400 30.400 ;
        RECT 86.000 29.800 88.400 30.400 ;
        RECT 82.800 29.600 83.600 29.800 ;
        RECT 79.600 28.800 80.200 29.600 ;
        RECT 79.200 28.200 80.200 28.800 ;
        RECT 79.200 28.000 80.000 28.200 ;
        RECT 81.200 27.600 82.000 29.200 ;
        RECT 84.400 27.600 85.200 29.200 ;
        RECT 77.600 27.400 78.400 27.600 ;
        RECT 77.600 27.000 80.600 27.400 ;
        RECT 77.600 26.800 81.800 27.000 ;
        RECT 80.000 26.400 81.800 26.800 ;
        RECT 81.200 26.200 81.800 26.400 ;
        RECT 86.000 26.200 86.600 29.800 ;
        RECT 87.600 29.600 88.400 29.800 ;
        RECT 90.800 28.800 91.600 30.400 ;
        RECT 92.200 28.400 92.800 31.800 ;
        RECT 94.000 31.700 96.400 31.800 ;
        RECT 94.000 31.600 94.800 31.700 ;
        RECT 95.600 31.600 96.400 31.700 ;
        RECT 97.600 28.400 98.200 31.800 ;
        RECT 102.800 30.400 103.600 30.800 ;
        RECT 106.800 30.400 107.400 31.800 ;
        RECT 98.800 28.800 99.600 30.400 ;
        RECT 102.000 29.800 103.600 30.400 ;
        RECT 105.200 29.800 107.600 30.400 ;
        RECT 102.000 29.600 102.800 29.800 ;
        RECT 89.200 28.200 90.000 28.400 ;
        RECT 89.200 27.600 90.800 28.200 ;
        RECT 92.200 27.600 94.800 28.400 ;
        RECT 95.600 27.600 98.200 28.400 ;
        RECT 100.400 28.300 101.200 28.400 ;
        RECT 102.100 28.300 102.700 29.600 ;
        RECT 100.400 28.200 102.700 28.300 ;
        RECT 99.600 27.700 102.700 28.200 ;
        RECT 99.600 27.600 101.200 27.700 ;
        RECT 103.600 27.600 104.400 29.200 ;
        RECT 90.000 27.200 90.800 27.600 ;
        RECT 76.400 25.200 77.800 26.200 ;
        RECT 77.000 22.200 77.800 25.200 ;
        RECT 81.200 22.200 82.000 26.200 ;
        RECT 86.000 22.200 86.800 26.200 ;
        RECT 87.600 25.600 88.400 26.400 ;
        RECT 89.400 26.200 93.000 26.600 ;
        RECT 94.000 26.200 94.600 27.600 ;
        RECT 95.800 26.200 96.400 27.600 ;
        RECT 99.600 27.200 100.400 27.600 ;
        RECT 97.400 26.200 101.000 26.600 ;
        RECT 105.200 26.200 105.800 29.800 ;
        RECT 106.800 29.600 107.600 29.800 ;
        RECT 108.400 28.300 109.200 39.800 ;
        RECT 114.200 32.400 115.000 39.800 ;
        RECT 115.600 33.600 116.400 34.400 ;
        RECT 115.800 32.400 116.400 33.600 ;
        RECT 120.600 32.400 121.400 39.800 ;
        RECT 122.000 33.600 122.800 34.400 ;
        RECT 122.200 32.400 122.800 33.600 ;
        RECT 125.000 32.600 125.800 39.800 ;
        RECT 114.200 31.800 115.200 32.400 ;
        RECT 115.800 31.800 117.200 32.400 ;
        RECT 120.600 31.800 121.600 32.400 ;
        RECT 122.200 31.800 123.600 32.400 ;
        RECT 125.000 31.800 126.800 32.600 ;
        RECT 113.200 28.800 114.000 30.400 ;
        RECT 114.600 28.400 115.200 31.800 ;
        RECT 116.400 31.600 117.200 31.800 ;
        RECT 119.600 28.800 120.400 30.400 ;
        RECT 121.000 30.300 121.600 31.800 ;
        RECT 122.800 31.600 123.600 31.800 ;
        RECT 124.400 30.300 125.200 31.200 ;
        RECT 121.000 29.700 125.200 30.300 ;
        RECT 121.000 28.400 121.600 29.700 ;
        RECT 124.400 29.600 125.200 29.700 ;
        RECT 126.000 30.300 126.600 31.800 ;
        RECT 134.000 31.400 134.800 39.800 ;
        RECT 138.400 36.400 139.200 39.800 ;
        RECT 137.200 35.800 139.200 36.400 ;
        RECT 142.800 35.800 143.600 39.800 ;
        RECT 147.000 35.800 148.200 39.800 ;
        RECT 137.200 35.000 138.000 35.800 ;
        RECT 142.800 35.200 143.400 35.800 ;
        RECT 140.600 34.600 144.200 35.200 ;
        RECT 146.800 35.000 147.600 35.800 ;
        RECT 140.600 34.400 141.400 34.600 ;
        RECT 143.400 34.400 144.200 34.600 ;
        RECT 137.200 33.000 138.000 33.200 ;
        RECT 141.800 33.000 142.600 33.200 ;
        RECT 137.200 32.400 142.600 33.000 ;
        RECT 143.200 33.000 145.400 33.600 ;
        RECT 143.200 31.800 143.800 33.000 ;
        RECT 144.600 32.800 145.400 33.000 ;
        RECT 147.000 33.200 148.400 34.000 ;
        RECT 147.000 32.200 147.600 33.200 ;
        RECT 139.000 31.400 143.800 31.800 ;
        RECT 134.000 31.200 143.800 31.400 ;
        RECT 145.200 31.600 147.600 32.200 ;
        RECT 134.000 31.000 139.800 31.200 ;
        RECT 134.000 30.800 139.600 31.000 ;
        RECT 132.400 30.300 133.200 30.400 ;
        RECT 126.000 29.700 133.200 30.300 ;
        RECT 140.400 30.200 141.200 30.400 ;
        RECT 126.000 28.400 126.600 29.700 ;
        RECT 132.400 29.600 133.200 29.700 ;
        RECT 136.200 29.600 141.200 30.200 ;
        RECT 136.200 29.400 137.000 29.600 ;
        RECT 138.800 29.400 139.600 29.600 ;
        RECT 137.800 28.400 138.600 28.600 ;
        RECT 145.200 28.400 145.800 31.600 ;
        RECT 151.600 31.200 152.400 39.800 ;
        RECT 148.200 30.600 152.400 31.200 ;
        RECT 148.200 30.400 149.000 30.600 ;
        RECT 149.800 29.800 150.600 30.000 ;
        RECT 146.800 29.200 150.600 29.800 ;
        RECT 146.800 29.000 147.600 29.200 ;
        RECT 111.600 28.300 112.400 28.400 ;
        RECT 108.400 28.200 112.400 28.300 ;
        RECT 108.400 27.700 113.200 28.200 ;
        RECT 89.200 26.000 93.200 26.200 ;
        RECT 87.400 24.800 88.200 25.600 ;
        RECT 89.200 22.200 90.000 26.000 ;
        RECT 92.400 22.200 93.200 26.000 ;
        RECT 94.000 22.200 94.800 26.200 ;
        RECT 95.600 22.200 96.400 26.200 ;
        RECT 97.200 26.000 101.200 26.200 ;
        RECT 97.200 22.200 98.000 26.000 ;
        RECT 100.400 22.200 101.200 26.000 ;
        RECT 105.200 22.200 106.000 26.200 ;
        RECT 106.800 25.600 107.600 26.400 ;
        RECT 106.600 24.800 107.400 25.600 ;
        RECT 108.400 22.200 109.200 27.700 ;
        RECT 111.600 27.600 113.200 27.700 ;
        RECT 114.600 27.600 117.200 28.400 ;
        RECT 118.000 28.200 118.800 28.400 ;
        RECT 118.000 27.600 119.600 28.200 ;
        RECT 121.000 27.600 123.600 28.400 ;
        RECT 126.000 27.600 126.800 28.400 ;
        RECT 134.800 27.800 145.800 28.400 ;
        RECT 134.800 27.600 136.400 27.800 ;
        RECT 112.400 27.200 113.200 27.600 ;
        RECT 110.000 24.800 110.800 26.400 ;
        RECT 111.800 26.200 115.400 26.600 ;
        RECT 116.400 26.200 117.000 27.600 ;
        RECT 118.800 27.200 119.600 27.600 ;
        RECT 118.200 26.200 121.800 26.600 ;
        RECT 122.800 26.200 123.400 27.600 ;
        RECT 111.600 26.000 115.600 26.200 ;
        RECT 111.600 22.200 112.400 26.000 ;
        RECT 114.800 22.200 115.600 26.000 ;
        RECT 116.400 22.200 117.200 26.200 ;
        RECT 118.000 26.000 122.000 26.200 ;
        RECT 118.000 22.200 118.800 26.000 ;
        RECT 121.200 22.200 122.000 26.000 ;
        RECT 122.800 22.200 123.600 26.200 ;
        RECT 126.000 24.200 126.600 27.600 ;
        RECT 126.000 22.200 126.800 24.200 ;
        RECT 134.000 22.200 134.800 27.000 ;
        RECT 139.000 25.600 139.600 27.800 ;
        RECT 142.000 27.600 142.800 27.800 ;
        RECT 144.600 27.600 145.400 27.800 ;
        RECT 151.600 27.200 152.400 30.600 ;
        RECT 148.600 26.600 152.400 27.200 ;
        RECT 148.600 26.400 149.400 26.600 ;
        RECT 137.200 24.200 138.000 25.000 ;
        RECT 138.800 24.800 139.600 25.600 ;
        RECT 140.600 25.400 141.400 25.600 ;
        RECT 140.600 24.800 143.400 25.400 ;
        RECT 142.800 24.200 143.400 24.800 ;
        RECT 146.800 24.200 147.600 25.000 ;
        RECT 137.200 23.600 139.200 24.200 ;
        RECT 138.400 22.200 139.200 23.600 ;
        RECT 142.800 22.200 143.600 24.200 ;
        RECT 146.800 23.600 148.200 24.200 ;
        RECT 147.000 22.200 148.200 23.600 ;
        RECT 151.600 22.200 152.400 26.600 ;
        RECT 153.200 31.200 154.000 39.800 ;
        RECT 157.400 35.800 158.600 39.800 ;
        RECT 162.000 35.800 162.800 39.800 ;
        RECT 166.400 36.400 167.200 39.800 ;
        RECT 166.400 35.800 168.400 36.400 ;
        RECT 158.000 35.000 158.800 35.800 ;
        RECT 162.200 35.200 162.800 35.800 ;
        RECT 161.400 34.600 165.000 35.200 ;
        RECT 167.600 35.000 168.400 35.800 ;
        RECT 161.400 34.400 162.200 34.600 ;
        RECT 164.200 34.400 165.000 34.600 ;
        RECT 157.200 33.200 158.600 34.000 ;
        RECT 158.000 32.200 158.600 33.200 ;
        RECT 160.200 33.000 162.400 33.600 ;
        RECT 160.200 32.800 161.000 33.000 ;
        RECT 158.000 31.600 160.400 32.200 ;
        RECT 153.200 30.600 157.400 31.200 ;
        RECT 153.200 27.200 154.000 30.600 ;
        RECT 156.600 30.400 157.400 30.600 ;
        RECT 159.800 30.400 160.400 31.600 ;
        RECT 161.800 31.800 162.400 33.000 ;
        RECT 163.000 33.000 163.800 33.200 ;
        RECT 167.600 33.000 168.400 33.200 ;
        RECT 163.000 32.400 168.400 33.000 ;
        RECT 161.800 31.400 166.600 31.800 ;
        RECT 170.800 31.400 171.600 39.800 ;
        RECT 161.800 31.200 171.600 31.400 ;
        RECT 165.800 31.000 171.600 31.200 ;
        RECT 166.000 30.800 171.600 31.000 ;
        RECT 172.400 31.400 173.200 39.800 ;
        RECT 176.800 36.400 177.600 39.800 ;
        RECT 175.600 35.800 177.600 36.400 ;
        RECT 181.200 35.800 182.000 39.800 ;
        RECT 185.400 35.800 186.600 39.800 ;
        RECT 175.600 35.000 176.400 35.800 ;
        RECT 181.200 35.200 181.800 35.800 ;
        RECT 179.000 34.600 182.600 35.200 ;
        RECT 185.200 35.000 186.000 35.800 ;
        RECT 179.000 34.400 179.800 34.600 ;
        RECT 181.800 34.400 182.600 34.600 ;
        RECT 175.600 33.000 176.400 33.200 ;
        RECT 180.200 33.000 181.000 33.200 ;
        RECT 175.600 32.400 181.000 33.000 ;
        RECT 181.600 33.000 183.800 33.600 ;
        RECT 181.600 31.800 182.200 33.000 ;
        RECT 183.000 32.800 183.800 33.000 ;
        RECT 185.400 33.200 186.800 34.000 ;
        RECT 185.400 32.200 186.000 33.200 ;
        RECT 177.400 31.400 182.200 31.800 ;
        RECT 172.400 31.200 182.200 31.400 ;
        RECT 183.600 31.600 186.000 32.200 ;
        RECT 172.400 31.000 178.200 31.200 ;
        RECT 172.400 30.800 178.000 31.000 ;
        RECT 155.000 29.800 155.800 30.000 ;
        RECT 155.000 29.200 158.800 29.800 ;
        RECT 159.600 29.600 160.400 30.400 ;
        RECT 164.400 30.200 165.200 30.400 ;
        RECT 178.800 30.200 179.600 30.400 ;
        RECT 164.400 29.600 169.400 30.200 ;
        RECT 158.000 29.000 158.800 29.200 ;
        RECT 159.800 28.400 160.400 29.600 ;
        RECT 166.000 29.400 166.800 29.600 ;
        RECT 168.600 29.400 169.400 29.600 ;
        RECT 174.600 29.600 179.600 30.200 ;
        RECT 174.600 29.400 175.400 29.600 ;
        RECT 167.000 28.400 167.800 28.600 ;
        RECT 176.200 28.400 177.000 28.600 ;
        RECT 183.600 28.400 184.200 31.600 ;
        RECT 190.000 31.200 190.800 39.800 ;
        RECT 186.600 30.600 190.800 31.200 ;
        RECT 186.600 30.400 187.400 30.600 ;
        RECT 188.200 29.800 189.000 30.000 ;
        RECT 185.200 29.200 189.000 29.800 ;
        RECT 185.200 29.000 186.000 29.200 ;
        RECT 159.800 28.300 170.800 28.400 ;
        RECT 173.200 28.300 184.200 28.400 ;
        RECT 159.800 27.800 184.200 28.300 ;
        RECT 160.200 27.600 161.000 27.800 ;
        RECT 153.200 26.600 157.200 27.200 ;
        RECT 153.200 22.200 154.000 26.600 ;
        RECT 156.200 26.400 157.200 26.600 ;
        RECT 156.400 26.300 157.200 26.400 ;
        RECT 159.600 26.300 160.400 26.400 ;
        RECT 156.400 25.700 160.400 26.300 ;
        RECT 159.600 25.600 160.400 25.700 ;
        RECT 166.000 25.600 166.600 27.800 ;
        RECT 169.200 27.700 174.800 27.800 ;
        RECT 169.200 27.600 170.800 27.700 ;
        RECT 173.200 27.600 174.800 27.700 ;
        RECT 164.200 25.400 165.000 25.600 ;
        RECT 158.000 24.200 158.800 25.000 ;
        RECT 162.200 24.800 165.000 25.400 ;
        RECT 166.000 24.800 166.800 25.600 ;
        RECT 162.200 24.200 162.800 24.800 ;
        RECT 167.600 24.200 168.400 25.000 ;
        RECT 157.400 23.600 158.800 24.200 ;
        RECT 157.400 22.200 158.600 23.600 ;
        RECT 162.000 22.200 162.800 24.200 ;
        RECT 166.400 23.600 168.400 24.200 ;
        RECT 166.400 22.200 167.200 23.600 ;
        RECT 170.800 22.200 171.600 27.000 ;
        RECT 172.400 22.200 173.200 27.000 ;
        RECT 177.400 25.600 178.000 27.800 ;
        RECT 183.000 27.600 183.800 27.800 ;
        RECT 190.000 27.200 190.800 30.600 ;
        RECT 187.000 26.600 190.800 27.200 ;
        RECT 187.000 26.400 187.800 26.600 ;
        RECT 175.600 24.200 176.400 25.000 ;
        RECT 177.200 24.800 178.000 25.600 ;
        RECT 179.000 25.400 179.800 25.600 ;
        RECT 179.000 24.800 181.800 25.400 ;
        RECT 181.200 24.200 181.800 24.800 ;
        RECT 185.200 24.200 186.000 25.000 ;
        RECT 175.600 23.600 177.600 24.200 ;
        RECT 176.800 22.200 177.600 23.600 ;
        RECT 181.200 22.200 182.000 24.200 ;
        RECT 185.200 23.600 186.600 24.200 ;
        RECT 185.400 22.200 186.600 23.600 ;
        RECT 190.000 22.200 190.800 26.600 ;
        RECT 4.400 15.200 5.200 19.800 ;
        RECT 3.000 14.600 5.200 15.200 ;
        RECT 6.000 15.400 6.800 19.800 ;
        RECT 10.200 18.400 11.400 19.800 ;
        RECT 10.200 17.800 11.600 18.400 ;
        RECT 14.800 17.800 15.600 19.800 ;
        RECT 19.200 18.400 20.000 19.800 ;
        RECT 19.200 17.800 21.200 18.400 ;
        RECT 10.800 17.000 11.600 17.800 ;
        RECT 15.000 17.200 15.600 17.800 ;
        RECT 15.000 16.600 17.800 17.200 ;
        RECT 17.000 16.400 17.800 16.600 ;
        RECT 18.800 16.400 19.600 17.200 ;
        RECT 20.400 17.000 21.200 17.800 ;
        RECT 9.000 15.400 9.800 15.600 ;
        RECT 6.000 14.800 9.800 15.400 ;
        RECT 3.000 11.600 3.600 14.600 ;
        RECT 4.400 11.600 5.200 13.200 ;
        RECT 2.400 10.800 3.600 11.600 ;
        RECT 3.000 10.200 3.600 10.800 ;
        RECT 6.000 11.400 6.800 14.800 ;
        RECT 13.000 14.200 13.800 14.400 ;
        RECT 17.200 14.200 18.000 14.400 ;
        RECT 18.800 14.200 19.400 16.400 ;
        RECT 23.600 15.000 24.400 19.800 ;
        RECT 25.400 16.400 26.200 17.200 ;
        RECT 25.200 15.600 26.000 16.400 ;
        RECT 26.800 15.800 27.600 19.800 ;
        RECT 32.200 16.800 33.000 19.800 ;
        RECT 22.000 14.200 23.600 14.400 ;
        RECT 12.600 13.600 23.600 14.200 ;
        RECT 10.800 12.800 11.600 13.000 ;
        RECT 7.800 12.200 11.600 12.800 ;
        RECT 7.800 12.000 8.600 12.200 ;
        RECT 9.400 11.400 10.200 11.600 ;
        RECT 6.000 10.800 10.200 11.400 ;
        RECT 3.000 9.600 5.200 10.200 ;
        RECT 4.400 2.200 5.200 9.600 ;
        RECT 6.000 2.200 6.800 10.800 ;
        RECT 12.600 10.400 13.200 13.600 ;
        RECT 19.800 13.400 20.600 13.600 ;
        RECT 18.800 12.400 19.600 12.600 ;
        RECT 21.400 12.400 22.200 12.600 ;
        RECT 17.200 11.800 22.200 12.400 ;
        RECT 25.200 12.200 26.000 12.400 ;
        RECT 27.000 12.200 27.600 15.800 ;
        RECT 31.600 15.800 33.000 16.800 ;
        RECT 36.400 15.800 37.200 19.800 ;
        RECT 41.200 15.800 42.000 19.800 ;
        RECT 46.000 17.800 46.800 19.800 ;
        RECT 42.600 16.400 43.400 17.200 ;
        RECT 42.800 16.300 43.600 16.400 ;
        RECT 44.400 16.300 45.200 16.400 ;
        RECT 28.400 12.800 29.200 14.400 ;
        RECT 31.600 12.400 32.200 15.800 ;
        RECT 36.400 15.600 37.000 15.800 ;
        RECT 35.200 15.200 37.000 15.600 ;
        RECT 32.800 15.000 37.000 15.200 ;
        RECT 32.800 14.600 35.800 15.000 ;
        RECT 32.800 14.400 33.600 14.600 ;
        RECT 30.000 12.200 30.800 12.400 ;
        RECT 17.200 11.600 18.000 11.800 ;
        RECT 25.200 11.600 27.600 12.200 ;
        RECT 29.200 11.600 30.800 12.200 ;
        RECT 31.600 11.600 32.400 12.400 ;
        RECT 18.800 11.000 24.400 11.200 ;
        RECT 18.600 10.800 24.400 11.000 ;
        RECT 10.800 9.800 13.200 10.400 ;
        RECT 14.600 10.600 24.400 10.800 ;
        RECT 14.600 10.200 19.400 10.600 ;
        RECT 10.800 8.800 11.400 9.800 ;
        RECT 10.000 8.000 11.400 8.800 ;
        RECT 13.000 9.000 13.800 9.200 ;
        RECT 14.600 9.000 15.200 10.200 ;
        RECT 13.000 8.400 15.200 9.000 ;
        RECT 15.800 9.000 21.200 9.600 ;
        RECT 15.800 8.800 16.600 9.000 ;
        RECT 20.400 8.800 21.200 9.000 ;
        RECT 14.200 7.400 15.000 7.600 ;
        RECT 17.000 7.400 17.800 7.600 ;
        RECT 10.800 6.200 11.600 7.000 ;
        RECT 14.200 6.800 17.800 7.400 ;
        RECT 15.000 6.200 15.600 6.800 ;
        RECT 20.400 6.200 21.200 7.000 ;
        RECT 10.200 2.200 11.400 6.200 ;
        RECT 14.800 2.200 15.600 6.200 ;
        RECT 19.200 5.600 21.200 6.200 ;
        RECT 19.200 2.200 20.000 5.600 ;
        RECT 23.600 2.200 24.400 10.600 ;
        RECT 25.400 10.200 26.000 11.600 ;
        RECT 29.200 11.200 30.000 11.600 ;
        RECT 31.600 10.200 32.200 11.600 ;
        RECT 33.000 11.000 33.600 14.400 ;
        RECT 36.400 12.800 37.200 14.400 ;
        RECT 39.600 12.800 40.400 14.400 ;
        RECT 38.000 12.200 38.800 12.400 ;
        RECT 41.200 12.200 41.800 15.800 ;
        RECT 42.800 15.700 45.200 16.300 ;
        RECT 42.800 15.600 43.600 15.700 ;
        RECT 44.400 15.600 45.200 15.700 ;
        RECT 46.000 14.400 46.600 17.800 ;
        RECT 47.600 15.600 48.400 17.200 ;
        RECT 54.000 15.000 54.800 19.800 ;
        RECT 58.400 18.400 59.200 19.800 ;
        RECT 57.200 17.800 59.200 18.400 ;
        RECT 62.800 17.800 63.600 19.800 ;
        RECT 67.000 18.400 68.200 19.800 ;
        RECT 66.800 17.800 68.200 18.400 ;
        RECT 57.200 17.000 58.000 17.800 ;
        RECT 62.800 17.200 63.400 17.800 ;
        RECT 58.800 16.400 59.600 17.200 ;
        RECT 60.600 16.600 63.400 17.200 ;
        RECT 66.800 17.000 67.600 17.800 ;
        RECT 60.600 16.400 61.400 16.600 ;
        RECT 46.000 13.600 46.800 14.400 ;
        RECT 54.800 14.200 56.400 14.400 ;
        RECT 59.000 14.200 59.600 16.400 ;
        RECT 68.600 15.400 69.400 15.600 ;
        RECT 71.600 15.400 72.400 19.800 ;
        RECT 68.600 14.800 72.400 15.400 ;
        RECT 76.400 15.200 77.200 19.800 ;
        RECT 64.600 14.200 65.400 14.400 ;
        RECT 54.800 13.600 65.800 14.200 ;
        RECT 42.800 12.300 43.600 12.400 ;
        RECT 44.400 12.300 45.200 12.400 ;
        RECT 42.800 12.200 45.200 12.300 ;
        RECT 38.000 11.600 39.600 12.200 ;
        RECT 41.200 11.700 45.200 12.200 ;
        RECT 41.200 11.600 43.600 11.700 ;
        RECT 38.800 11.200 39.600 11.600 ;
        RECT 33.000 10.400 35.400 11.000 ;
        RECT 25.200 2.200 26.000 10.200 ;
        RECT 26.800 9.600 30.800 10.200 ;
        RECT 26.800 2.200 27.600 9.600 ;
        RECT 30.000 2.200 30.800 9.600 ;
        RECT 31.600 2.200 32.400 10.200 ;
        RECT 34.800 6.200 35.400 10.400 ;
        RECT 42.800 10.200 43.400 11.600 ;
        RECT 44.400 10.800 45.200 11.700 ;
        RECT 46.000 12.300 46.600 13.600 ;
        RECT 57.800 13.400 58.600 13.600 ;
        RECT 56.200 12.400 57.000 12.600 ;
        RECT 58.800 12.400 59.600 12.600 ;
        RECT 52.400 12.300 53.200 12.400 ;
        RECT 46.000 11.700 53.200 12.300 ;
        RECT 56.200 11.800 61.200 12.400 ;
        RECT 46.000 10.200 46.600 11.700 ;
        RECT 52.400 11.600 53.200 11.700 ;
        RECT 60.400 11.600 61.200 11.800 ;
        RECT 54.000 11.000 59.600 11.200 ;
        RECT 54.000 10.800 59.800 11.000 ;
        RECT 54.000 10.600 63.800 10.800 ;
        RECT 38.000 9.600 42.000 10.200 ;
        RECT 34.800 2.200 35.600 6.200 ;
        RECT 38.000 2.200 38.800 9.600 ;
        RECT 41.200 2.200 42.000 9.600 ;
        RECT 42.800 2.200 43.600 10.200 ;
        RECT 45.000 9.400 46.800 10.200 ;
        RECT 45.000 2.200 45.800 9.400 ;
        RECT 54.000 2.200 54.800 10.600 ;
        RECT 59.000 10.200 63.800 10.600 ;
        RECT 57.200 9.000 62.600 9.600 ;
        RECT 57.200 8.800 58.000 9.000 ;
        RECT 61.800 8.800 62.600 9.000 ;
        RECT 63.200 9.000 63.800 10.200 ;
        RECT 65.200 10.400 65.800 13.600 ;
        RECT 66.800 12.800 67.600 13.000 ;
        RECT 66.800 12.200 70.600 12.800 ;
        RECT 69.800 12.000 70.600 12.200 ;
        RECT 68.200 11.400 69.000 11.600 ;
        RECT 71.600 11.400 72.400 14.800 ;
        RECT 75.000 14.600 77.200 15.200 ;
        RECT 78.000 15.200 78.800 19.800 ;
        RECT 82.800 15.200 83.600 19.800 ;
        RECT 87.600 15.200 88.400 19.800 ;
        RECT 92.400 15.200 93.200 19.800 ;
        RECT 97.200 15.400 98.000 19.800 ;
        RECT 101.400 18.400 102.600 19.800 ;
        RECT 101.400 17.800 102.800 18.400 ;
        RECT 106.000 17.800 106.800 19.800 ;
        RECT 110.400 18.400 111.200 19.800 ;
        RECT 110.400 17.800 112.400 18.400 ;
        RECT 102.000 17.000 102.800 17.800 ;
        RECT 106.200 17.200 106.800 17.800 ;
        RECT 106.200 16.600 109.000 17.200 ;
        RECT 108.200 16.400 109.000 16.600 ;
        RECT 110.000 16.400 110.800 17.200 ;
        RECT 111.600 17.000 112.400 17.800 ;
        RECT 100.200 15.400 101.000 15.600 ;
        RECT 78.000 14.600 80.200 15.200 ;
        RECT 82.800 14.600 85.000 15.200 ;
        RECT 87.600 14.600 89.800 15.200 ;
        RECT 92.400 14.600 94.600 15.200 ;
        RECT 75.000 11.600 75.600 14.600 ;
        RECT 76.400 11.600 77.200 13.200 ;
        RECT 78.000 11.600 78.800 13.200 ;
        RECT 79.600 11.600 80.200 14.600 ;
        RECT 82.800 11.600 83.600 13.200 ;
        RECT 84.400 11.600 85.000 14.600 ;
        RECT 87.600 11.600 88.400 13.200 ;
        RECT 89.200 11.600 89.800 14.600 ;
        RECT 92.400 11.600 93.200 13.200 ;
        RECT 94.000 11.600 94.600 14.600 ;
        RECT 97.200 14.800 101.000 15.400 ;
        RECT 68.200 10.800 72.400 11.400 ;
        RECT 74.400 10.800 75.600 11.600 ;
        RECT 65.200 9.800 67.600 10.400 ;
        RECT 64.600 9.000 65.400 9.200 ;
        RECT 63.200 8.400 65.400 9.000 ;
        RECT 67.000 8.800 67.600 9.800 ;
        RECT 67.000 8.000 68.400 8.800 ;
        RECT 60.600 7.400 61.400 7.600 ;
        RECT 63.400 7.400 64.200 7.600 ;
        RECT 57.200 6.200 58.000 7.000 ;
        RECT 60.600 6.800 64.200 7.400 ;
        RECT 62.800 6.200 63.400 6.800 ;
        RECT 66.800 6.200 67.600 7.000 ;
        RECT 57.200 5.600 59.200 6.200 ;
        RECT 58.400 2.200 59.200 5.600 ;
        RECT 62.800 2.200 63.600 6.200 ;
        RECT 67.000 2.200 68.200 6.200 ;
        RECT 71.600 2.200 72.400 10.800 ;
        RECT 75.000 10.200 75.600 10.800 ;
        RECT 79.600 10.800 80.800 11.600 ;
        RECT 84.400 10.800 85.600 11.600 ;
        RECT 89.200 10.800 90.400 11.600 ;
        RECT 94.000 10.800 95.200 11.600 ;
        RECT 97.200 11.400 98.000 14.800 ;
        RECT 104.200 14.200 105.000 14.400 ;
        RECT 106.800 14.200 107.600 14.400 ;
        RECT 110.000 14.200 110.600 16.400 ;
        RECT 114.800 15.000 115.600 19.800 ;
        RECT 117.000 18.400 117.800 19.800 ;
        RECT 117.000 17.600 118.800 18.400 ;
        RECT 117.000 16.400 117.800 17.600 ;
        RECT 117.000 15.800 118.800 16.400 ;
        RECT 113.200 14.200 114.800 14.400 ;
        RECT 103.800 13.600 114.800 14.200 ;
        RECT 102.000 12.800 102.800 13.000 ;
        RECT 99.000 12.200 102.800 12.800 ;
        RECT 99.000 12.000 99.800 12.200 ;
        RECT 100.600 11.400 101.400 11.600 ;
        RECT 97.200 10.800 101.400 11.400 ;
        RECT 79.600 10.200 80.200 10.800 ;
        RECT 84.400 10.200 85.000 10.800 ;
        RECT 89.200 10.200 89.800 10.800 ;
        RECT 94.000 10.200 94.600 10.800 ;
        RECT 75.000 9.600 77.200 10.200 ;
        RECT 76.400 2.200 77.200 9.600 ;
        RECT 78.000 9.600 80.200 10.200 ;
        RECT 82.800 9.600 85.000 10.200 ;
        RECT 87.600 9.600 89.800 10.200 ;
        RECT 92.400 9.600 94.600 10.200 ;
        RECT 78.000 2.200 78.800 9.600 ;
        RECT 82.800 2.200 83.600 9.600 ;
        RECT 87.600 2.200 88.400 9.600 ;
        RECT 92.400 2.200 93.200 9.600 ;
        RECT 97.200 2.200 98.000 10.800 ;
        RECT 103.800 10.400 104.400 13.600 ;
        RECT 111.000 13.400 111.800 13.600 ;
        RECT 112.600 12.400 113.400 12.600 ;
        RECT 108.400 11.800 113.400 12.400 ;
        RECT 108.400 11.600 109.200 11.800 ;
        RECT 110.000 11.000 115.600 11.200 ;
        RECT 109.800 10.800 115.600 11.000 ;
        RECT 102.000 9.800 104.400 10.400 ;
        RECT 105.800 10.600 115.600 10.800 ;
        RECT 105.800 10.200 110.600 10.600 ;
        RECT 102.000 8.800 102.600 9.800 ;
        RECT 101.200 8.000 102.600 8.800 ;
        RECT 104.200 9.000 105.000 9.200 ;
        RECT 105.800 9.000 106.400 10.200 ;
        RECT 104.200 8.400 106.400 9.000 ;
        RECT 107.000 9.000 112.400 9.600 ;
        RECT 107.000 8.800 107.800 9.000 ;
        RECT 111.600 8.800 112.400 9.000 ;
        RECT 105.400 7.400 106.200 7.600 ;
        RECT 108.200 7.400 109.000 7.600 ;
        RECT 102.000 6.200 102.800 7.000 ;
        RECT 105.400 6.800 109.000 7.400 ;
        RECT 106.200 6.200 106.800 6.800 ;
        RECT 111.600 6.200 112.400 7.000 ;
        RECT 101.400 2.200 102.600 6.200 ;
        RECT 106.000 2.200 106.800 6.200 ;
        RECT 110.400 5.600 112.400 6.200 ;
        RECT 110.400 2.200 111.200 5.600 ;
        RECT 114.800 2.200 115.600 10.600 ;
        RECT 116.400 8.800 117.200 10.400 ;
        RECT 118.000 2.200 118.800 15.800 ;
        RECT 119.600 13.600 120.400 15.200 ;
        RECT 121.200 15.000 122.000 19.800 ;
        RECT 125.600 18.400 126.400 19.800 ;
        RECT 124.400 17.800 126.400 18.400 ;
        RECT 130.000 17.800 130.800 19.800 ;
        RECT 134.200 18.400 135.400 19.800 ;
        RECT 134.000 17.800 135.400 18.400 ;
        RECT 124.400 17.000 125.200 17.800 ;
        RECT 130.000 17.200 130.600 17.800 ;
        RECT 126.000 16.400 126.800 17.200 ;
        RECT 127.800 16.600 130.600 17.200 ;
        RECT 134.000 17.000 134.800 17.800 ;
        RECT 127.800 16.400 128.600 16.600 ;
        RECT 122.000 14.200 123.600 14.400 ;
        RECT 126.200 14.200 126.800 16.400 ;
        RECT 135.800 15.400 136.600 15.600 ;
        RECT 138.800 15.400 139.600 19.800 ;
        RECT 135.800 14.800 139.600 15.400 ;
        RECT 131.800 14.200 132.600 14.400 ;
        RECT 122.000 13.600 133.000 14.200 ;
        RECT 125.000 13.400 125.800 13.600 ;
        RECT 123.400 12.400 124.200 12.600 ;
        RECT 126.000 12.400 126.800 12.600 ;
        RECT 123.400 11.800 128.400 12.400 ;
        RECT 127.600 11.600 128.400 11.800 ;
        RECT 121.200 11.000 126.800 11.200 ;
        RECT 121.200 10.800 127.000 11.000 ;
        RECT 121.200 10.600 131.000 10.800 ;
        RECT 121.200 2.200 122.000 10.600 ;
        RECT 126.200 10.200 131.000 10.600 ;
        RECT 124.400 9.000 129.800 9.600 ;
        RECT 124.400 8.800 125.200 9.000 ;
        RECT 129.000 8.800 129.800 9.000 ;
        RECT 130.400 9.000 131.000 10.200 ;
        RECT 132.400 10.400 133.000 13.600 ;
        RECT 134.000 12.800 134.800 13.000 ;
        RECT 134.000 12.200 137.800 12.800 ;
        RECT 137.000 12.000 137.800 12.200 ;
        RECT 138.800 12.300 139.600 14.800 ;
        RECT 145.200 15.200 146.000 19.800 ;
        RECT 150.000 15.200 150.800 19.800 ;
        RECT 154.800 15.200 155.600 19.800 ;
        RECT 159.600 15.200 160.400 19.800 ;
        RECT 164.400 15.600 165.200 17.200 ;
        RECT 145.200 14.600 147.400 15.200 ;
        RECT 150.000 14.600 152.200 15.200 ;
        RECT 154.800 14.600 157.000 15.200 ;
        RECT 159.600 14.600 161.800 15.200 ;
        RECT 145.200 12.300 146.000 13.200 ;
        RECT 138.800 11.700 146.000 12.300 ;
        RECT 135.400 11.400 136.200 11.600 ;
        RECT 138.800 11.400 139.600 11.700 ;
        RECT 145.200 11.600 146.000 11.700 ;
        RECT 146.800 11.600 147.400 14.600 ;
        RECT 150.000 11.600 150.800 13.200 ;
        RECT 151.600 11.600 152.200 14.600 ;
        RECT 154.800 11.600 155.600 13.200 ;
        RECT 156.400 11.600 157.000 14.600 ;
        RECT 159.600 11.600 160.400 13.200 ;
        RECT 161.200 11.600 161.800 14.600 ;
        RECT 166.000 14.300 166.800 19.800 ;
        RECT 170.800 15.800 171.600 19.800 ;
        RECT 175.600 17.800 176.400 19.800 ;
        RECT 169.200 14.300 170.000 14.400 ;
        RECT 166.000 13.700 170.000 14.300 ;
        RECT 135.400 10.800 139.600 11.400 ;
        RECT 132.400 9.800 134.800 10.400 ;
        RECT 131.800 9.000 132.600 9.200 ;
        RECT 130.400 8.400 132.600 9.000 ;
        RECT 134.200 8.800 134.800 9.800 ;
        RECT 134.200 8.000 135.600 8.800 ;
        RECT 127.800 7.400 128.600 7.600 ;
        RECT 130.600 7.400 131.400 7.600 ;
        RECT 124.400 6.200 125.200 7.000 ;
        RECT 127.800 6.800 131.400 7.400 ;
        RECT 130.000 6.200 130.600 6.800 ;
        RECT 134.000 6.200 134.800 7.000 ;
        RECT 124.400 5.600 126.400 6.200 ;
        RECT 125.600 2.200 126.400 5.600 ;
        RECT 130.000 2.200 130.800 6.200 ;
        RECT 134.200 2.200 135.400 6.200 ;
        RECT 138.800 2.200 139.600 10.800 ;
        RECT 146.800 10.800 148.000 11.600 ;
        RECT 151.600 10.800 152.800 11.600 ;
        RECT 156.400 10.800 157.600 11.600 ;
        RECT 161.200 10.800 162.400 11.600 ;
        RECT 146.800 10.200 147.400 10.800 ;
        RECT 151.600 10.200 152.200 10.800 ;
        RECT 156.400 10.200 157.000 10.800 ;
        RECT 161.200 10.200 161.800 10.800 ;
        RECT 145.200 9.600 147.400 10.200 ;
        RECT 150.000 9.600 152.200 10.200 ;
        RECT 154.800 9.600 157.000 10.200 ;
        RECT 159.600 9.600 161.800 10.200 ;
        RECT 145.200 2.200 146.000 9.600 ;
        RECT 150.000 2.200 150.800 9.600 ;
        RECT 154.800 2.200 155.600 9.600 ;
        RECT 159.600 2.200 160.400 9.600 ;
        RECT 166.000 2.200 166.800 13.700 ;
        RECT 169.200 12.800 170.000 13.700 ;
        RECT 167.600 12.200 168.400 12.400 ;
        RECT 170.800 12.200 171.400 15.800 ;
        RECT 174.000 15.600 174.800 17.200 ;
        RECT 175.800 15.600 176.400 17.800 ;
        RECT 178.800 15.800 179.600 19.800 ;
        RECT 181.000 18.400 181.800 19.800 ;
        RECT 180.400 17.600 181.800 18.400 ;
        RECT 181.000 16.800 181.800 17.600 ;
        RECT 175.800 15.000 178.200 15.600 ;
        RECT 175.600 13.600 176.600 14.400 ;
        RECT 176.000 12.800 176.800 13.600 ;
        RECT 172.400 12.200 173.200 12.400 ;
        RECT 167.600 11.600 169.200 12.200 ;
        RECT 170.800 11.600 173.200 12.200 ;
        RECT 177.600 12.000 178.200 15.000 ;
        RECT 179.000 14.400 179.600 15.800 ;
        RECT 178.800 13.600 179.600 14.400 ;
        RECT 179.000 12.400 179.600 13.600 ;
        RECT 168.400 11.200 169.200 11.600 ;
        RECT 172.400 10.200 173.000 11.600 ;
        RECT 177.400 11.400 178.200 12.000 ;
        RECT 178.800 11.600 179.600 12.400 ;
        RECT 174.000 11.200 178.200 11.400 ;
        RECT 174.000 10.800 178.000 11.200 ;
        RECT 167.600 9.600 171.600 10.200 ;
        RECT 167.600 2.200 168.400 9.600 ;
        RECT 170.800 2.200 171.600 9.600 ;
        RECT 172.400 2.200 173.200 10.200 ;
        RECT 174.000 2.200 174.800 10.800 ;
        RECT 179.000 10.200 179.600 11.600 ;
        RECT 178.200 9.600 179.600 10.200 ;
        RECT 180.400 15.800 181.800 16.800 ;
        RECT 185.200 15.800 186.000 19.800 ;
        RECT 187.000 16.400 187.800 17.200 ;
        RECT 180.400 12.400 181.000 15.800 ;
        RECT 185.200 15.600 185.800 15.800 ;
        RECT 186.800 15.600 187.600 16.400 ;
        RECT 188.400 15.800 189.200 19.800 ;
        RECT 184.000 15.200 185.800 15.600 ;
        RECT 181.600 15.000 185.800 15.200 ;
        RECT 181.600 14.600 184.600 15.000 ;
        RECT 181.600 14.400 182.400 14.600 ;
        RECT 180.400 11.600 181.200 12.400 ;
        RECT 180.400 10.200 181.000 11.600 ;
        RECT 181.800 11.000 182.400 14.400 ;
        RECT 183.200 13.800 184.000 14.000 ;
        RECT 183.200 13.200 184.200 13.800 ;
        RECT 183.600 12.400 184.200 13.200 ;
        RECT 185.200 12.800 186.000 14.400 ;
        RECT 183.600 11.600 184.400 12.400 ;
        RECT 186.800 12.200 187.600 12.400 ;
        RECT 188.600 12.200 189.200 15.800 ;
        RECT 190.000 12.800 190.800 14.400 ;
        RECT 191.600 12.200 192.400 12.400 ;
        RECT 186.800 11.600 189.200 12.200 ;
        RECT 190.800 11.600 192.400 12.200 ;
        RECT 181.800 10.400 184.200 11.000 ;
        RECT 178.200 2.200 179.000 9.600 ;
        RECT 180.400 2.200 181.200 10.200 ;
        RECT 183.600 6.200 184.200 10.400 ;
        RECT 187.000 10.200 187.600 11.600 ;
        RECT 190.800 11.200 191.600 11.600 ;
        RECT 183.600 2.200 184.400 6.200 ;
        RECT 186.800 2.200 187.600 10.200 ;
        RECT 188.400 9.600 192.400 10.200 ;
        RECT 188.400 2.200 189.200 9.600 ;
        RECT 191.600 2.200 192.400 9.600 ;
      LAYER via1 ;
        RECT 26.800 173.600 27.600 174.400 ;
        RECT 20.400 172.200 21.200 173.000 ;
        RECT 12.400 163.600 13.200 164.400 ;
        RECT 28.400 171.800 29.200 172.600 ;
        RECT 41.200 173.600 42.000 174.400 ;
        RECT 33.200 170.200 34.000 171.000 ;
        RECT 15.600 163.600 16.400 164.400 ;
        RECT 39.600 170.200 40.400 171.000 ;
        RECT 94.000 173.600 94.800 174.400 ;
        RECT 82.800 172.200 83.600 173.000 ;
        RECT 90.800 171.800 91.600 172.600 ;
        RECT 95.600 170.200 96.400 171.000 ;
        RECT 78.000 163.600 78.800 164.400 ;
        RECT 111.600 172.200 112.400 173.000 ;
        RECT 119.600 171.800 120.400 172.600 ;
        RECT 124.400 170.200 125.200 171.000 ;
        RECT 182.000 177.600 182.800 178.400 ;
        RECT 145.200 172.200 146.000 173.000 ;
        RECT 153.200 171.800 154.000 172.600 ;
        RECT 166.000 173.600 166.800 174.400 ;
        RECT 106.800 163.600 107.600 164.400 ;
        RECT 158.000 170.200 158.800 171.000 ;
        RECT 140.400 167.600 141.200 168.400 ;
        RECT 164.400 170.200 165.200 171.000 ;
        RECT 15.600 152.400 16.400 153.200 ;
        RECT 18.800 151.000 19.600 151.800 ;
        RECT 34.800 152.400 35.600 153.200 ;
        RECT 38.000 151.000 38.800 151.800 ;
        RECT 39.600 157.600 40.400 158.400 ;
        RECT 18.800 146.200 19.600 147.000 ;
        RECT 1.200 143.600 2.000 144.400 ;
        RECT 38.000 146.200 38.800 147.000 ;
        RECT 20.400 143.600 21.200 144.400 ;
        RECT 42.800 148.000 43.600 148.800 ;
        RECT 46.000 145.600 46.800 146.400 ;
        RECT 65.200 145.600 66.000 146.400 ;
        RECT 63.600 143.600 64.400 144.400 ;
        RECT 78.000 147.600 78.800 148.400 ;
        RECT 81.200 147.600 82.000 148.400 ;
        RECT 100.400 157.600 101.200 158.400 ;
        RECT 86.000 147.600 86.800 148.400 ;
        RECT 87.600 145.600 88.400 146.400 ;
        RECT 113.200 157.600 114.000 158.400 ;
        RECT 126.000 149.600 126.800 150.400 ;
        RECT 129.200 147.600 130.000 148.400 ;
        RECT 156.400 153.600 157.200 154.400 ;
        RECT 146.800 149.600 147.600 150.400 ;
        RECT 159.600 151.600 160.400 152.400 ;
        RECT 170.800 152.400 171.600 153.200 ;
        RECT 174.000 151.000 174.800 151.800 ;
        RECT 154.800 145.600 155.600 146.400 ;
        RECT 174.000 146.200 174.800 147.000 ;
        RECT 175.600 146.200 176.400 147.000 ;
        RECT 193.200 143.600 194.000 144.400 ;
        RECT 14.000 137.600 14.800 138.400 ;
        RECT 12.400 133.600 13.200 134.400 ;
        RECT 25.200 135.600 26.000 136.400 ;
        RECT 20.400 133.600 21.200 134.400 ;
        RECT 22.000 129.600 22.800 130.400 ;
        RECT 31.600 137.600 32.400 138.400 ;
        RECT 28.400 133.600 29.200 134.400 ;
        RECT 41.200 137.600 42.000 138.400 ;
        RECT 34.800 133.600 35.600 134.400 ;
        RECT 30.000 129.600 30.800 130.400 ;
        RECT 44.400 131.600 45.200 132.400 ;
        RECT 46.000 125.600 46.800 126.400 ;
        RECT 65.200 137.600 66.000 138.400 ;
        RECT 68.400 137.600 69.200 138.400 ;
        RECT 58.800 133.600 59.600 134.400 ;
        RECT 49.200 123.600 50.000 124.400 ;
        RECT 63.600 129.600 64.400 130.400 ;
        RECT 84.400 137.600 85.200 138.400 ;
        RECT 79.600 129.600 80.400 130.400 ;
        RECT 103.600 137.600 104.400 138.400 ;
        RECT 100.400 133.600 101.200 134.400 ;
        RECT 89.200 132.200 90.000 133.000 ;
        RECT 108.400 132.200 109.200 133.000 ;
        RECT 102.000 130.200 102.800 131.000 ;
        RECT 121.200 130.200 122.000 131.000 ;
        RECT 126.000 131.600 126.800 132.400 ;
        RECT 127.600 129.600 128.400 130.400 ;
        RECT 145.200 135.600 146.000 136.400 ;
        RECT 135.600 133.600 136.400 134.400 ;
        RECT 137.200 131.600 138.000 132.400 ;
        RECT 129.200 123.600 130.000 124.400 ;
        RECT 154.800 137.600 155.600 138.400 ;
        RECT 153.200 133.600 154.000 134.400 ;
        RECT 150.000 131.600 150.800 132.400 ;
        RECT 170.800 137.600 171.600 138.400 ;
        RECT 161.200 133.600 162.000 134.400 ;
        RECT 162.800 129.600 163.600 130.400 ;
        RECT 172.400 133.600 173.200 134.400 ;
        RECT 177.200 133.600 178.000 134.400 ;
        RECT 167.600 129.600 168.400 130.400 ;
        RECT 174.000 131.600 174.800 132.400 ;
        RECT 175.600 130.200 176.400 131.000 ;
        RECT 193.200 123.600 194.000 124.400 ;
        RECT 6.000 113.600 6.800 114.400 ;
        RECT 4.400 109.600 5.200 110.400 ;
        RECT 20.400 112.400 21.200 113.200 ;
        RECT 23.600 111.000 24.400 111.800 ;
        RECT 23.600 106.200 24.400 107.000 ;
        RECT 46.000 117.600 46.800 118.400 ;
        RECT 60.400 117.600 61.200 118.400 ;
        RECT 47.600 113.600 48.400 114.400 ;
        RECT 58.800 113.600 59.600 114.400 ;
        RECT 41.200 109.600 42.000 110.400 ;
        RECT 50.800 111.600 51.600 112.400 ;
        RECT 49.200 109.600 50.000 110.400 ;
        RECT 60.400 109.600 61.200 110.400 ;
        RECT 34.800 105.600 35.600 106.400 ;
        RECT 70.000 107.600 70.800 108.400 ;
        RECT 74.800 105.600 75.600 106.400 ;
        RECT 79.600 107.600 80.400 108.400 ;
        RECT 87.600 109.600 88.400 110.400 ;
        RECT 86.000 107.600 86.800 108.400 ;
        RECT 89.200 107.600 90.000 108.400 ;
        RECT 76.400 103.600 77.200 104.400 ;
        RECT 82.800 103.600 83.600 104.400 ;
        RECT 114.800 112.400 115.600 113.200 ;
        RECT 138.800 113.600 139.600 114.400 ;
        RECT 118.000 111.000 118.800 111.800 ;
        RECT 166.000 117.600 166.800 118.400 ;
        RECT 172.400 113.600 173.200 114.400 ;
        RECT 185.200 117.600 186.000 118.400 ;
        RECT 98.800 105.600 99.600 106.400 ;
        RECT 126.000 107.600 126.800 108.400 ;
        RECT 118.000 106.200 118.800 107.000 ;
        RECT 122.800 105.600 123.600 106.400 ;
        RECT 124.400 106.200 125.200 107.000 ;
        RECT 121.200 103.600 122.000 104.400 ;
        RECT 156.400 109.600 157.200 110.400 ;
        RECT 169.200 111.600 170.000 112.400 ;
        RECT 167.600 105.600 168.400 106.400 ;
        RECT 188.400 109.600 189.200 110.400 ;
        RECT 17.200 93.600 18.000 94.400 ;
        RECT 49.200 97.600 50.000 98.400 ;
        RECT 10.800 92.200 11.600 93.000 ;
        RECT 18.800 91.800 19.600 92.600 ;
        RECT 23.600 90.200 24.400 91.000 ;
        RECT 6.000 83.600 6.800 84.400 ;
        RECT 30.000 89.600 30.800 90.400 ;
        RECT 36.400 91.600 37.200 92.400 ;
        RECT 63.600 97.600 64.400 98.400 ;
        RECT 47.600 89.600 48.400 90.400 ;
        RECT 58.800 93.600 59.600 94.400 ;
        RECT 74.800 97.600 75.600 98.400 ;
        RECT 68.400 89.600 69.200 90.400 ;
        RECT 89.200 97.600 90.000 98.400 ;
        RECT 79.600 91.600 80.400 92.400 ;
        RECT 111.600 97.600 112.400 98.400 ;
        RECT 94.000 92.200 94.800 93.000 ;
        RECT 106.800 90.200 107.600 91.000 ;
        RECT 122.800 97.600 123.600 98.400 ;
        RECT 121.200 93.600 122.000 94.400 ;
        RECT 134.000 93.600 134.800 94.400 ;
        RECT 129.200 91.600 130.000 92.400 ;
        RECT 130.800 91.600 131.600 92.400 ;
        RECT 145.200 93.600 146.000 94.400 ;
        RECT 148.400 93.600 149.200 94.400 ;
        RECT 156.400 93.600 157.200 94.400 ;
        RECT 158.000 91.600 158.800 92.400 ;
        RECT 153.200 83.600 154.000 84.400 ;
        RECT 180.400 83.600 181.200 84.400 ;
        RECT 9.200 77.600 10.000 78.400 ;
        RECT 7.600 73.600 8.400 74.400 ;
        RECT 4.400 69.600 5.200 70.400 ;
        RECT 10.800 71.600 11.600 72.400 ;
        RECT 9.200 69.600 10.000 70.400 ;
        RECT 14.000 69.600 14.800 70.400 ;
        RECT 23.600 67.600 24.400 68.400 ;
        RECT 22.000 65.600 22.800 66.400 ;
        RECT 30.000 77.600 30.800 78.400 ;
        RECT 33.200 69.600 34.000 70.400 ;
        RECT 60.400 73.600 61.200 74.400 ;
        RECT 30.000 67.600 30.800 68.400 ;
        RECT 41.200 65.600 42.000 66.400 ;
        RECT 42.800 66.200 43.600 67.000 ;
        RECT 47.600 65.600 48.400 66.400 ;
        RECT 68.400 77.600 69.200 78.400 ;
        RECT 86.000 77.600 86.800 78.400 ;
        RECT 73.200 69.600 74.000 70.400 ;
        RECT 89.200 69.600 90.000 70.400 ;
        RECT 70.000 63.600 70.800 64.400 ;
        RECT 97.200 69.600 98.000 70.400 ;
        RECT 95.600 67.600 96.400 68.400 ;
        RECT 98.800 67.600 99.600 68.400 ;
        RECT 108.400 67.600 109.200 68.400 ;
        RECT 106.800 66.200 107.600 67.000 ;
        RECT 127.600 69.600 128.400 70.400 ;
        RECT 130.800 69.600 131.600 70.400 ;
        RECT 126.000 65.600 126.800 66.400 ;
        RECT 146.800 71.600 147.600 72.400 ;
        RECT 150.000 67.600 150.800 68.400 ;
        RECT 169.200 72.400 170.000 73.200 ;
        RECT 172.400 71.000 173.200 71.800 ;
        RECT 191.600 77.600 192.400 78.400 ;
        RECT 175.600 67.600 176.400 68.400 ;
        RECT 167.600 65.600 168.400 66.400 ;
        RECT 153.200 63.600 154.000 64.400 ;
        RECT 154.800 63.600 155.600 64.400 ;
        RECT 172.400 66.200 173.200 67.000 ;
        RECT 174.000 66.200 174.800 67.000 ;
        RECT 6.000 57.600 6.800 58.400 ;
        RECT 17.200 53.600 18.000 54.400 ;
        RECT 30.000 57.600 30.800 58.400 ;
        RECT 22.000 53.600 22.800 54.400 ;
        RECT 10.800 52.200 11.600 53.000 ;
        RECT 18.800 51.800 19.600 52.600 ;
        RECT 23.600 50.200 24.400 51.000 ;
        RECT 31.600 53.600 32.400 54.400 ;
        RECT 52.400 53.600 53.200 54.400 ;
        RECT 50.800 50.200 51.600 51.000 ;
        RECT 68.400 43.600 69.200 44.400 ;
        RECT 73.200 49.600 74.000 50.400 ;
        RECT 89.200 55.600 90.000 56.400 ;
        RECT 82.800 53.600 83.600 54.400 ;
        RECT 84.400 51.600 85.200 52.400 ;
        RECT 89.200 49.600 90.000 50.400 ;
        RECT 105.200 49.600 106.000 50.400 ;
        RECT 102.000 43.600 102.800 44.400 ;
        RECT 122.800 57.600 123.600 58.400 ;
        RECT 121.200 51.600 122.000 52.400 ;
        RECT 132.400 49.600 133.200 50.400 ;
        RECT 143.600 53.600 144.400 54.400 ;
        RECT 145.200 49.600 146.000 50.400 ;
        RECT 150.000 53.600 150.800 54.400 ;
        RECT 164.400 57.600 165.200 58.400 ;
        RECT 154.800 49.600 155.600 50.400 ;
        RECT 166.000 51.600 166.800 52.400 ;
        RECT 172.400 51.600 173.200 52.400 ;
        RECT 161.200 43.600 162.000 44.400 ;
        RECT 15.600 32.400 16.400 33.200 ;
        RECT 18.800 31.000 19.600 31.800 ;
        RECT 23.600 29.600 24.400 30.400 ;
        RECT 18.800 26.200 19.600 27.000 ;
        RECT 25.200 27.600 26.000 28.400 ;
        RECT 1.200 23.600 2.000 24.400 ;
        RECT 20.400 23.600 21.200 24.400 ;
        RECT 26.800 25.600 27.600 26.400 ;
        RECT 36.400 27.600 37.200 28.400 ;
        RECT 46.000 29.600 46.800 30.400 ;
        RECT 68.400 33.600 69.200 34.400 ;
        RECT 73.200 37.600 74.000 38.400 ;
        RECT 71.600 33.600 72.400 34.400 ;
        RECT 47.600 27.600 48.400 28.400 ;
        RECT 42.800 23.600 43.600 24.400 ;
        RECT 73.200 29.600 74.000 30.400 ;
        RECT 90.800 29.600 91.600 30.400 ;
        RECT 98.800 29.600 99.600 30.400 ;
        RECT 92.400 27.600 93.200 28.400 ;
        RECT 97.200 27.600 98.000 28.400 ;
        RECT 108.400 29.600 109.200 30.400 ;
        RECT 113.200 29.600 114.000 30.400 ;
        RECT 119.600 29.600 120.400 30.400 ;
        RECT 86.000 23.600 86.800 24.400 ;
        RECT 105.200 23.600 106.000 24.400 ;
        RECT 116.400 27.600 117.200 28.400 ;
        RECT 110.000 25.600 110.800 26.400 ;
        RECT 134.000 26.200 134.800 27.000 ;
        RECT 151.600 23.600 152.400 24.400 ;
        RECT 153.200 37.600 154.000 38.400 ;
        RECT 167.600 32.400 168.400 33.200 ;
        RECT 170.800 31.000 171.600 31.800 ;
        RECT 190.000 37.600 190.800 38.400 ;
        RECT 178.800 29.600 179.600 30.400 ;
        RECT 170.800 26.200 171.600 27.000 ;
        RECT 172.400 26.200 173.200 27.000 ;
        RECT 6.000 17.600 6.800 18.400 ;
        RECT 17.200 13.600 18.000 14.400 ;
        RECT 10.800 12.200 11.600 13.000 ;
        RECT 18.800 11.800 19.600 12.600 ;
        RECT 28.400 13.600 29.200 14.400 ;
        RECT 23.600 10.200 24.400 11.000 ;
        RECT 30.000 11.600 30.800 12.400 ;
        RECT 36.400 13.600 37.200 14.400 ;
        RECT 39.600 13.600 40.400 14.400 ;
        RECT 71.600 17.600 72.400 18.400 ;
        RECT 55.600 13.600 56.400 14.400 ;
        RECT 58.800 11.800 59.600 12.600 ;
        RECT 54.000 10.200 54.800 11.000 ;
        RECT 97.200 17.600 98.000 18.400 ;
        RECT 106.800 13.600 107.600 14.400 ;
        RECT 118.000 17.600 118.800 18.400 ;
        RECT 102.000 12.200 102.800 13.000 ;
        RECT 114.800 10.200 115.600 11.000 ;
        RECT 116.400 9.600 117.200 10.400 ;
        RECT 138.800 17.600 139.600 18.400 ;
        RECT 122.800 13.600 123.600 14.400 ;
        RECT 126.000 11.800 126.800 12.600 ;
        RECT 121.200 10.200 122.000 11.000 ;
        RECT 169.200 13.600 170.000 14.400 ;
        RECT 172.400 11.600 173.200 12.400 ;
        RECT 188.400 17.600 189.200 18.400 ;
        RECT 185.200 13.600 186.000 14.400 ;
        RECT 190.000 13.600 190.800 14.400 ;
        RECT 191.600 11.600 192.400 12.400 ;
      LAYER metal2 ;
        RECT 20.400 166.200 21.200 177.800 ;
        RECT 26.800 173.600 27.600 174.400 ;
        RECT 12.400 163.600 13.200 164.400 ;
        RECT 15.600 163.600 16.400 164.400 ;
        RECT 1.200 143.600 2.000 144.400 ;
        RECT 6.000 144.200 6.800 155.800 ;
        RECT 12.500 150.400 13.100 163.600 ;
        RECT 15.700 160.400 16.300 163.600 ;
        RECT 15.600 159.600 16.400 160.400 ;
        RECT 23.600 159.600 24.400 160.400 ;
        RECT 12.400 149.600 13.200 150.400 ;
        RECT 12.500 148.400 13.100 149.600 ;
        RECT 14.000 149.400 14.800 150.200 ;
        RECT 12.400 147.600 13.200 148.400 ;
        RECT 9.200 143.600 10.000 144.400 ;
        RECT 1.300 132.400 1.900 143.600 ;
        RECT 9.300 132.400 9.900 143.600 ;
        RECT 14.100 138.400 14.700 149.400 ;
        RECT 15.600 144.200 16.400 155.800 ;
        RECT 17.200 147.600 18.000 148.400 ;
        RECT 14.000 137.600 14.800 138.400 ;
        RECT 15.600 135.600 16.400 136.400 ;
        RECT 12.400 133.600 13.200 134.400 ;
        RECT 15.600 133.600 16.400 134.400 ;
        RECT 1.200 131.600 2.000 132.400 ;
        RECT 4.400 131.600 5.200 132.400 ;
        RECT 9.200 131.600 10.000 132.400 ;
        RECT 10.800 131.600 11.600 132.400 ;
        RECT 12.500 130.400 13.100 133.600 ;
        RECT 15.700 132.400 16.300 133.600 ;
        RECT 15.600 131.600 16.400 132.400 ;
        RECT 12.400 129.600 13.200 130.400 ;
        RECT 6.000 113.600 6.800 114.400 ;
        RECT 6.100 110.400 6.700 113.600 ;
        RECT 4.400 109.600 5.200 110.400 ;
        RECT 6.000 109.600 6.800 110.400 ;
        RECT 10.800 104.200 11.600 115.800 ;
        RECT 17.300 108.400 17.900 147.600 ;
        RECT 18.800 146.200 19.600 151.800 ;
        RECT 20.400 143.600 21.200 144.400 ;
        RECT 23.700 136.400 24.300 159.600 ;
        RECT 25.200 144.200 26.000 155.800 ;
        RECT 26.900 150.400 27.500 173.600 ;
        RECT 28.400 171.800 29.200 172.600 ;
        RECT 28.500 166.400 29.100 171.800 ;
        RECT 28.400 165.600 29.200 166.400 ;
        RECT 30.000 166.200 30.800 177.800 ;
        RECT 33.200 170.200 34.000 175.800 ;
        RECT 34.800 171.600 35.600 172.400 ;
        RECT 34.900 160.400 35.500 171.600 ;
        RECT 39.600 170.200 40.400 175.800 ;
        RECT 41.200 173.600 42.000 174.400 ;
        RECT 39.600 165.600 40.400 166.400 ;
        RECT 42.800 166.200 43.600 177.800 ;
        RECT 46.000 171.600 46.800 172.400 ;
        RECT 46.100 166.400 46.700 171.600 ;
        RECT 46.000 165.600 46.800 166.400 ;
        RECT 52.400 166.200 53.200 177.800 ;
        RECT 63.600 171.600 64.400 172.400 ;
        RECT 68.400 171.600 69.200 172.400 ;
        RECT 73.200 171.600 74.000 172.400 ;
        RECT 34.800 159.600 35.600 160.400 ;
        RECT 39.700 158.400 40.300 165.600 ;
        RECT 58.800 163.600 59.600 164.400 ;
        RECT 39.600 157.600 40.400 158.400 ;
        RECT 26.800 149.600 27.600 150.400 ;
        RECT 33.200 149.400 34.000 150.400 ;
        RECT 31.600 145.600 32.400 146.400 ;
        RECT 30.000 143.600 30.800 144.400 ;
        RECT 20.400 135.600 21.200 136.400 ;
        RECT 23.600 135.600 24.400 136.400 ;
        RECT 25.200 135.600 26.000 136.400 ;
        RECT 20.500 134.400 21.100 135.600 ;
        RECT 23.700 134.400 24.300 135.600 ;
        RECT 20.400 133.600 21.200 134.400 ;
        RECT 23.600 133.600 24.400 134.400 ;
        RECT 26.800 133.600 27.600 134.400 ;
        RECT 28.400 133.600 29.200 134.400 ;
        RECT 18.800 131.600 19.600 132.400 ;
        RECT 18.900 130.400 19.500 131.600 ;
        RECT 30.100 130.400 30.700 143.600 ;
        RECT 31.700 138.400 32.300 145.600 ;
        RECT 34.800 144.200 35.600 155.800 ;
        RECT 58.900 152.400 59.500 163.600 ;
        RECT 63.700 152.400 64.300 171.600 ;
        RECT 68.500 152.400 69.100 171.600 ;
        RECT 73.300 166.400 73.900 171.600 ;
        RECT 70.000 165.600 70.800 166.400 ;
        RECT 73.200 165.600 74.000 166.400 ;
        RECT 78.000 165.600 78.800 166.400 ;
        RECT 82.800 166.200 83.600 177.800 ;
        RECT 90.800 171.800 91.600 172.600 ;
        RECT 90.900 170.400 91.500 171.800 ;
        RECT 90.800 169.600 91.600 170.400 ;
        RECT 92.400 166.200 93.200 177.800 ;
        RECT 94.000 173.600 94.800 174.400 ;
        RECT 95.600 170.200 96.400 175.800 ;
        RECT 100.400 171.600 101.200 172.400 ;
        RECT 105.200 171.600 106.000 172.400 ;
        RECT 100.400 169.600 101.200 170.400 ;
        RECT 38.000 146.200 38.800 151.800 ;
        RECT 58.800 151.600 59.600 152.400 ;
        RECT 63.600 152.300 64.400 152.400 ;
        RECT 62.100 151.700 64.400 152.300 ;
        RECT 49.200 149.600 50.000 150.400 ;
        RECT 52.400 149.600 53.200 150.400 ;
        RECT 42.800 148.300 43.600 148.800 ;
        RECT 41.300 148.000 43.600 148.300 ;
        RECT 41.300 147.700 43.500 148.000 ;
        RECT 41.300 138.400 41.900 147.700 ;
        RECT 44.400 147.600 45.200 148.400 ;
        RECT 44.500 146.400 45.100 147.600 ;
        RECT 49.300 146.400 49.900 149.600 ;
        RECT 58.800 147.600 59.600 148.400 ;
        RECT 44.400 145.600 45.200 146.400 ;
        RECT 46.000 145.600 46.800 146.400 ;
        RECT 49.200 145.600 50.000 146.400 ;
        RECT 54.000 145.600 54.800 146.400 ;
        RECT 46.100 144.400 46.700 145.600 ;
        RECT 54.100 144.400 54.700 145.600 ;
        RECT 46.000 143.600 46.800 144.400 ;
        RECT 54.000 143.600 54.800 144.400 ;
        RECT 31.600 137.600 32.400 138.400 ;
        RECT 41.200 137.600 42.000 138.400 ;
        RECT 34.800 135.600 35.600 136.400 ;
        RECT 36.400 136.300 37.200 136.400 ;
        RECT 36.400 135.700 38.700 136.300 ;
        RECT 36.400 135.600 37.200 135.700 ;
        RECT 34.900 134.400 35.500 135.600 ;
        RECT 34.800 133.600 35.600 134.400 ;
        RECT 38.100 132.400 38.700 135.700 ;
        RECT 47.600 135.600 48.400 136.400 ;
        RECT 50.800 135.600 51.600 136.400 ;
        RECT 58.900 134.400 59.500 147.600 ;
        RECT 62.100 138.400 62.700 151.700 ;
        RECT 63.600 151.600 64.400 151.700 ;
        RECT 65.200 151.600 66.000 152.400 ;
        RECT 68.400 151.600 69.200 152.400 ;
        RECT 65.300 146.400 65.900 151.600 ;
        RECT 70.100 150.400 70.700 165.600 ;
        RECT 78.100 164.400 78.700 165.600 ;
        RECT 78.000 163.600 78.800 164.400 ;
        RECT 74.800 151.600 75.600 152.400 ;
        RECT 70.000 149.600 70.800 150.400 ;
        RECT 73.200 149.600 74.000 150.400 ;
        RECT 78.100 148.400 78.700 163.600 ;
        RECT 100.500 158.400 101.100 169.600 ;
        RECT 100.400 157.600 101.200 158.400 ;
        RECT 95.600 151.600 96.400 152.400 ;
        RECT 82.800 149.600 83.600 150.400 ;
        RECT 89.200 150.300 90.000 150.400 ;
        RECT 87.700 149.700 90.000 150.300 ;
        RECT 68.400 147.600 69.200 148.400 ;
        RECT 71.600 147.600 72.400 148.400 ;
        RECT 78.000 147.600 78.800 148.400 ;
        RECT 81.200 147.600 82.000 148.400 ;
        RECT 86.000 147.600 86.800 148.400 ;
        RECT 87.700 146.400 88.300 149.700 ;
        RECT 89.200 149.600 90.000 149.700 ;
        RECT 94.000 149.600 94.800 150.400 ;
        RECT 95.700 150.300 96.300 151.600 ;
        RECT 97.200 150.300 98.000 150.400 ;
        RECT 95.700 149.700 98.000 150.300 ;
        RECT 97.200 149.600 98.000 149.700 ;
        RECT 94.100 148.400 94.700 149.600 ;
        RECT 94.000 147.600 94.800 148.400 ;
        RECT 65.200 145.600 66.000 146.400 ;
        RECT 68.400 145.600 69.200 146.400 ;
        RECT 87.600 145.600 88.400 146.400 ;
        RECT 63.600 143.600 64.400 144.400 ;
        RECT 65.200 143.600 66.000 144.400 ;
        RECT 62.000 137.600 62.800 138.400 ;
        RECT 62.100 136.400 62.700 137.600 ;
        RECT 63.700 136.400 64.300 143.600 ;
        RECT 65.300 138.400 65.900 143.600 ;
        RECT 68.500 138.400 69.100 145.600 ;
        RECT 74.800 143.600 75.600 144.400 ;
        RECT 65.200 137.600 66.000 138.400 ;
        RECT 68.400 137.600 69.200 138.400 ;
        RECT 62.000 135.600 62.800 136.400 ;
        RECT 63.600 135.600 64.400 136.400 ;
        RECT 74.900 134.400 75.500 143.600 ;
        RECT 84.400 137.600 85.200 138.400 ;
        RECT 44.400 133.600 45.200 134.400 ;
        RECT 58.800 133.600 59.600 134.400 ;
        RECT 66.800 133.600 67.600 134.400 ;
        RECT 74.800 133.600 75.600 134.400 ;
        RECT 82.800 134.300 83.600 134.400 ;
        RECT 82.800 133.700 85.100 134.300 ;
        RECT 82.800 133.600 83.600 133.700 ;
        RECT 44.500 132.400 45.100 133.600 ;
        RECT 58.900 132.400 59.500 133.600 ;
        RECT 38.000 131.600 38.800 132.400 ;
        RECT 44.400 131.600 45.200 132.400 ;
        RECT 57.200 131.600 58.000 132.400 ;
        RECT 58.800 131.600 59.600 132.400 ;
        RECT 63.600 131.600 64.400 132.400 ;
        RECT 18.800 129.600 19.600 130.400 ;
        RECT 22.000 129.600 22.800 130.400 ;
        RECT 30.000 129.600 30.800 130.400 ;
        RECT 36.400 129.600 37.200 130.400 ;
        RECT 18.800 111.600 19.600 112.400 ;
        RECT 18.900 110.200 19.500 111.600 ;
        RECT 18.800 109.400 19.600 110.200 ;
        RECT 17.200 107.600 18.000 108.400 ;
        RECT 9.200 91.600 10.000 92.400 ;
        RECT 6.000 84.300 6.800 84.400 ;
        RECT 6.000 83.700 8.300 84.300 ;
        RECT 6.000 83.600 6.800 83.700 ;
        RECT 7.700 74.400 8.300 83.700 ;
        RECT 9.300 78.400 9.900 91.600 ;
        RECT 10.800 86.200 11.600 97.800 ;
        RECT 12.400 95.600 13.200 96.400 ;
        RECT 17.300 94.400 17.900 107.600 ;
        RECT 20.400 104.200 21.200 115.800 ;
        RECT 22.100 108.400 22.700 129.600 ;
        RECT 36.500 128.400 37.100 129.600 ;
        RECT 36.400 127.600 37.200 128.400 ;
        RECT 36.500 118.400 37.100 127.600 ;
        RECT 38.100 124.400 38.700 131.600 ;
        RECT 57.300 128.400 57.900 131.600 ;
        RECT 63.600 129.600 64.400 130.400 ;
        RECT 66.900 130.300 67.500 133.600 ;
        RECT 71.600 131.600 72.400 132.400 ;
        RECT 73.200 131.600 74.000 132.400 ;
        RECT 68.400 130.300 69.200 130.400 ;
        RECT 66.900 129.700 69.200 130.300 ;
        RECT 68.400 129.600 69.200 129.700 ;
        RECT 63.700 128.400 64.300 129.600 ;
        RECT 71.700 128.400 72.300 131.600 ;
        RECT 57.200 127.600 58.000 128.400 ;
        RECT 60.400 127.600 61.200 128.400 ;
        RECT 63.600 127.600 64.400 128.400 ;
        RECT 71.600 127.600 72.400 128.400 ;
        RECT 46.000 125.600 46.800 126.400 ;
        RECT 38.000 123.600 38.800 124.400 ;
        RECT 46.000 123.600 46.800 124.400 ;
        RECT 49.200 123.600 50.000 124.400 ;
        RECT 46.100 118.400 46.700 123.600 ;
        RECT 36.400 117.600 37.200 118.400 ;
        RECT 41.200 117.600 42.000 118.400 ;
        RECT 46.000 117.600 46.800 118.400 ;
        RECT 38.000 113.600 38.800 114.400 ;
        RECT 47.600 113.600 48.400 114.400 ;
        RECT 22.000 107.600 22.800 108.400 ;
        RECT 23.600 106.200 24.400 111.800 ;
        RECT 25.200 111.600 26.000 112.400 ;
        RECT 28.400 109.600 29.200 110.400 ;
        RECT 30.000 107.600 30.800 108.400 ;
        RECT 17.200 93.600 18.000 94.400 ;
        RECT 18.800 93.600 19.600 94.400 ;
        RECT 18.900 92.600 19.500 93.600 ;
        RECT 18.800 91.800 19.600 92.600 ;
        RECT 20.400 86.200 21.200 97.800 ;
        RECT 23.600 90.200 24.400 95.800 ;
        RECT 25.200 95.600 26.000 96.400 ;
        RECT 25.300 94.400 25.900 95.600 ;
        RECT 25.200 93.600 26.000 94.400 ;
        RECT 26.800 91.600 27.600 92.400 ;
        RECT 26.900 82.400 27.500 91.600 ;
        RECT 30.100 90.400 30.700 107.600 ;
        RECT 34.800 105.600 35.600 106.400 ;
        RECT 38.100 98.400 38.700 113.600 ;
        RECT 44.400 111.600 45.200 112.400 ;
        RECT 47.600 111.600 48.400 112.400 ;
        RECT 41.200 109.600 42.000 110.400 ;
        RECT 39.600 107.600 40.400 108.400 ;
        RECT 39.700 106.400 40.300 107.600 ;
        RECT 39.600 105.600 40.400 106.400 ;
        RECT 38.000 97.600 38.800 98.400 ;
        RECT 39.700 96.400 40.300 105.600 ;
        RECT 41.300 98.400 41.900 109.600 ;
        RECT 44.500 108.400 45.100 111.600 ;
        RECT 44.400 107.600 45.200 108.400 ;
        RECT 41.200 97.600 42.000 98.400 ;
        RECT 46.000 97.600 46.800 98.400 ;
        RECT 39.600 95.600 40.400 96.400 ;
        RECT 41.200 95.600 42.000 96.400 ;
        RECT 31.600 93.600 32.400 94.400 ;
        RECT 41.300 92.400 41.900 95.600 ;
        RECT 36.400 91.600 37.200 92.400 ;
        RECT 41.200 91.600 42.000 92.400 ;
        RECT 44.400 91.600 45.200 92.400 ;
        RECT 47.700 90.400 48.300 111.600 ;
        RECT 49.300 110.400 49.900 123.600 ;
        RECT 60.500 118.400 61.100 127.600 ;
        RECT 65.200 125.600 66.000 126.400 ;
        RECT 60.400 117.600 61.200 118.400 ;
        RECT 58.800 113.600 59.600 114.400 ;
        RECT 50.800 111.600 51.600 112.400 ;
        RECT 63.600 111.600 64.400 112.400 ;
        RECT 49.200 109.600 50.000 110.400 ;
        RECT 60.400 109.600 61.200 110.400 ;
        RECT 63.700 108.400 64.300 111.600 ;
        RECT 65.300 110.400 65.900 125.600 ;
        RECT 70.000 111.600 70.800 112.400 ;
        RECT 73.200 111.600 74.000 112.400 ;
        RECT 65.200 109.600 66.000 110.400 ;
        RECT 73.200 109.600 74.000 110.400 ;
        RECT 49.200 107.600 50.000 108.400 ;
        RECT 63.600 107.600 64.400 108.400 ;
        RECT 70.000 107.600 70.800 108.400 ;
        RECT 49.300 98.400 49.900 107.600 ;
        RECT 63.700 102.400 64.300 107.600 ;
        RECT 63.600 101.600 64.400 102.400 ;
        RECT 49.200 97.600 50.000 98.400 ;
        RECT 63.600 97.600 64.400 98.400 ;
        RECT 68.400 97.600 69.200 98.400 ;
        RECT 63.700 96.400 64.300 97.600 ;
        RECT 63.600 95.600 64.400 96.400 ;
        RECT 58.800 93.600 59.600 94.400 ;
        RECT 54.000 91.600 54.800 92.400 ;
        RECT 60.400 91.600 61.200 92.400 ;
        RECT 54.100 90.400 54.700 91.600 ;
        RECT 68.500 90.400 69.100 97.600 ;
        RECT 70.100 96.400 70.700 107.600 ;
        RECT 74.900 106.400 75.500 133.600 ;
        RECT 79.600 131.600 80.400 132.400 ;
        RECT 84.500 130.400 85.100 133.700 ;
        RECT 79.600 129.600 80.400 130.400 ;
        RECT 84.400 129.600 85.200 130.400 ;
        RECT 78.000 127.600 78.800 128.400 ;
        RECT 78.100 110.400 78.700 127.600 ;
        RECT 79.700 124.400 80.300 129.600 ;
        RECT 79.600 123.600 80.400 124.400 ;
        RECT 84.500 112.400 85.100 129.600 ;
        RECT 87.700 128.400 88.300 145.600 ;
        RECT 87.600 127.600 88.400 128.400 ;
        RECT 89.200 126.200 90.000 137.800 ;
        RECT 95.600 131.600 96.400 132.400 ;
        RECT 98.800 126.200 99.600 137.800 ;
        RECT 103.600 137.600 104.400 138.400 ;
        RECT 100.400 133.600 101.200 134.400 ;
        RECT 102.000 130.200 102.800 135.800 ;
        RECT 103.700 130.400 104.300 137.600 ;
        RECT 105.300 134.400 105.900 171.600 ;
        RECT 111.600 166.200 112.400 177.800 ;
        RECT 113.200 173.600 114.000 174.400 ;
        RECT 113.300 172.400 113.900 173.600 ;
        RECT 113.200 171.600 114.000 172.400 ;
        RECT 119.600 171.800 120.400 172.600 ;
        RECT 106.800 163.600 107.600 164.400 ;
        RECT 106.900 148.400 107.500 163.600 ;
        RECT 113.300 158.400 113.900 171.600 ;
        RECT 113.200 157.600 114.000 158.400 ;
        RECT 119.700 150.400 120.300 171.800 ;
        RECT 121.200 166.200 122.000 177.800 ;
        RECT 124.400 170.200 125.200 175.800 ;
        RECT 126.000 171.600 126.800 172.400 ;
        RECT 130.800 171.600 131.600 172.400 ;
        RECT 126.100 160.400 126.700 171.600 ;
        RECT 130.900 168.400 131.500 171.600 ;
        RECT 130.800 167.600 131.600 168.400 ;
        RECT 140.400 167.600 141.200 168.400 ;
        RECT 126.000 159.600 126.800 160.400 ;
        RECT 129.200 159.600 130.000 160.400 ;
        RECT 122.800 151.600 123.600 152.400 ;
        RECT 116.400 149.600 117.200 150.400 ;
        RECT 118.000 149.600 118.800 150.400 ;
        RECT 119.600 149.600 120.400 150.400 ;
        RECT 126.000 149.600 126.800 150.400 ;
        RECT 116.500 148.400 117.100 149.600 ;
        RECT 118.100 148.400 118.700 149.600 ;
        RECT 129.300 148.400 129.900 159.600 ;
        RECT 106.800 147.600 107.600 148.400 ;
        RECT 116.400 147.600 117.200 148.400 ;
        RECT 118.000 147.600 118.800 148.400 ;
        RECT 129.200 147.600 130.000 148.400 ;
        RECT 118.100 146.300 118.700 147.600 ;
        RECT 116.500 145.700 118.700 146.300 ;
        RECT 105.200 133.600 106.000 134.400 ;
        RECT 103.600 129.600 104.400 130.400 ;
        RECT 108.400 126.200 109.200 137.800 ;
        RECT 110.000 133.600 110.800 134.400 ;
        RECT 110.100 132.400 110.700 133.600 ;
        RECT 110.000 131.600 110.800 132.400 ;
        RECT 114.800 131.600 115.600 132.400 ;
        RECT 98.800 123.600 99.600 124.400 ;
        RECT 98.900 114.400 99.500 123.600 ;
        RECT 98.800 113.600 99.600 114.400 ;
        RECT 82.800 111.600 83.600 112.400 ;
        RECT 84.400 111.600 85.200 112.400 ;
        RECT 92.400 111.600 93.200 112.400 ;
        RECT 82.900 110.400 83.500 111.600 ;
        RECT 78.000 109.600 78.800 110.400 ;
        RECT 82.800 109.600 83.600 110.400 ;
        RECT 79.600 107.600 80.400 108.400 ;
        RECT 74.800 106.300 75.600 106.400 ;
        RECT 73.300 105.700 75.600 106.300 ;
        RECT 73.300 96.400 73.900 105.700 ;
        RECT 74.800 105.600 75.600 105.700 ;
        RECT 79.700 104.400 80.300 107.600 ;
        RECT 84.500 104.400 85.100 111.600 ;
        RECT 92.500 110.400 93.100 111.600 ;
        RECT 87.600 109.600 88.400 110.400 ;
        RECT 92.400 109.600 93.200 110.400 ;
        RECT 94.000 109.600 94.800 110.400 ;
        RECT 94.100 108.400 94.700 109.600 ;
        RECT 86.000 107.600 86.800 108.400 ;
        RECT 89.200 107.600 90.000 108.400 ;
        RECT 94.000 107.600 94.800 108.400 ;
        RECT 95.600 107.600 96.400 108.400 ;
        RECT 86.100 106.400 86.700 107.600 ;
        RECT 98.900 106.400 99.500 113.600 ;
        RECT 86.000 105.600 86.800 106.400 ;
        RECT 90.800 105.600 91.600 106.400 ;
        RECT 98.800 105.600 99.600 106.400 ;
        RECT 74.800 103.600 75.600 104.400 ;
        RECT 76.400 103.600 77.200 104.400 ;
        RECT 79.600 103.600 80.400 104.400 ;
        RECT 82.800 103.600 83.600 104.400 ;
        RECT 84.400 103.600 85.200 104.400 ;
        RECT 105.200 104.200 106.000 115.800 ;
        RECT 110.100 110.400 110.700 131.600 ;
        RECT 111.600 111.600 112.400 112.400 ;
        RECT 111.700 110.400 112.300 111.600 ;
        RECT 110.000 109.600 110.800 110.400 ;
        RECT 111.600 109.600 112.400 110.400 ;
        RECT 110.100 108.400 110.700 109.600 ;
        RECT 110.000 107.600 110.800 108.400 ;
        RECT 111.600 107.600 112.400 108.400 ;
        RECT 74.900 98.400 75.500 103.600 ;
        RECT 74.800 97.600 75.600 98.400 ;
        RECT 70.000 95.600 70.800 96.400 ;
        RECT 73.200 95.600 74.000 96.400 ;
        RECT 70.000 93.600 70.800 94.400 ;
        RECT 76.500 92.400 77.100 103.600 ;
        RECT 82.900 96.400 83.500 103.600 ;
        RECT 84.400 97.600 85.200 98.400 ;
        RECT 89.200 97.600 90.000 98.400 ;
        RECT 84.500 96.400 85.100 97.600 ;
        RECT 82.800 95.600 83.600 96.400 ;
        RECT 84.400 95.600 85.200 96.400 ;
        RECT 87.600 95.600 88.400 96.400 ;
        RECT 76.400 91.600 77.200 92.400 ;
        RECT 78.000 91.600 78.800 92.400 ;
        RECT 79.600 91.600 80.400 92.400 ;
        RECT 87.600 91.600 88.400 92.400 ;
        RECT 78.100 90.400 78.700 91.600 ;
        RECT 30.000 89.600 30.800 90.400 ;
        RECT 47.600 89.600 48.400 90.400 ;
        RECT 54.000 89.600 54.800 90.400 ;
        RECT 68.400 89.600 69.200 90.400 ;
        RECT 73.200 89.600 74.000 90.400 ;
        RECT 78.000 89.600 78.800 90.400 ;
        RECT 89.200 89.600 90.000 90.400 ;
        RECT 30.100 84.400 30.700 89.600 ;
        RECT 30.000 83.600 30.800 84.400 ;
        RECT 36.400 83.600 37.200 84.400 ;
        RECT 26.800 81.600 27.600 82.400 ;
        RECT 30.000 81.600 30.800 82.400 ;
        RECT 30.100 78.400 30.700 81.600 ;
        RECT 9.200 77.600 10.000 78.400 ;
        RECT 30.000 77.600 30.800 78.400 ;
        RECT 7.600 73.600 8.400 74.400 ;
        RECT 36.500 72.400 37.100 83.600 ;
        RECT 73.300 78.400 73.900 89.600 ;
        RECT 86.000 81.600 86.800 82.400 ;
        RECT 86.100 78.400 86.700 81.600 ;
        RECT 68.400 77.600 69.200 78.400 ;
        RECT 73.200 77.600 74.000 78.400 ;
        RECT 86.000 77.600 86.800 78.400 ;
        RECT 10.800 71.600 11.600 72.400 ;
        RECT 14.000 71.600 14.800 72.400 ;
        RECT 17.200 71.600 18.000 72.400 ;
        RECT 26.800 71.600 27.600 72.400 ;
        RECT 36.400 71.600 37.200 72.400 ;
        RECT 39.600 71.600 40.400 72.400 ;
        RECT 14.100 70.400 14.700 71.600 ;
        RECT 4.400 69.600 5.200 70.400 ;
        RECT 9.200 69.600 10.000 70.400 ;
        RECT 14.000 69.600 14.800 70.400 ;
        RECT 23.600 69.600 24.400 70.400 ;
        RECT 14.100 58.400 14.700 69.600 ;
        RECT 23.700 68.400 24.300 69.600 ;
        RECT 23.600 67.600 24.400 68.400 ;
        RECT 26.900 66.400 27.500 71.600 ;
        RECT 31.600 69.600 32.400 70.400 ;
        RECT 33.200 69.600 34.000 70.400 ;
        RECT 38.000 69.600 38.800 70.400 ;
        RECT 31.700 68.400 32.300 69.600 ;
        RECT 30.000 67.600 30.800 68.400 ;
        RECT 31.600 67.600 32.400 68.400 ;
        RECT 33.300 66.400 33.900 69.600 ;
        RECT 38.100 68.400 38.700 69.600 ;
        RECT 38.000 67.600 38.800 68.400 ;
        RECT 18.800 65.600 19.600 66.400 ;
        RECT 22.000 65.600 22.800 66.400 ;
        RECT 26.800 65.600 27.600 66.400 ;
        RECT 30.000 65.600 30.800 66.400 ;
        RECT 33.200 65.600 34.000 66.400 ;
        RECT 38.000 65.600 38.800 66.400 ;
        RECT 41.200 65.600 42.000 66.400 ;
        RECT 42.800 66.200 43.600 71.800 ;
        RECT 6.000 57.600 6.800 58.400 ;
        RECT 10.800 46.200 11.600 57.800 ;
        RECT 14.000 57.600 14.800 58.400 ;
        RECT 17.200 53.600 18.000 54.400 ;
        RECT 1.200 23.600 2.000 24.400 ;
        RECT 4.400 23.600 5.200 24.400 ;
        RECT 6.000 24.200 6.800 35.800 ;
        RECT 14.000 29.400 14.800 30.400 ;
        RECT 15.600 24.200 16.400 35.800 ;
        RECT 17.300 28.400 17.900 53.600 ;
        RECT 18.900 52.600 19.500 65.600 ;
        RECT 30.100 58.400 30.700 65.600 ;
        RECT 46.000 64.200 46.800 75.800 ;
        RECT 47.600 71.600 48.400 72.400 ;
        RECT 47.700 70.200 48.300 71.600 ;
        RECT 47.600 69.400 48.400 70.200 ;
        RECT 47.600 65.600 48.400 66.400 ;
        RECT 18.800 51.800 19.600 52.600 ;
        RECT 20.400 46.200 21.200 57.800 ;
        RECT 26.800 57.600 27.600 58.400 ;
        RECT 30.000 57.600 30.800 58.400 ;
        RECT 22.000 53.600 22.800 54.400 ;
        RECT 23.600 50.200 24.400 55.800 ;
        RECT 26.900 54.000 27.500 57.600 ;
        RECT 47.700 54.400 48.300 65.600 ;
        RECT 55.600 64.200 56.400 75.800 ;
        RECT 60.400 73.600 61.200 74.400 ;
        RECT 60.500 70.400 61.100 73.600 ;
        RECT 73.300 70.400 73.900 77.600 ;
        RECT 89.300 70.400 89.900 89.600 ;
        RECT 94.000 86.200 94.800 97.800 ;
        RECT 95.600 91.600 96.400 92.400 ;
        RECT 98.800 91.600 99.600 92.400 ;
        RECT 95.700 82.400 96.300 91.600 ;
        RECT 103.600 86.200 104.400 97.800 ;
        RECT 106.800 90.200 107.600 95.800 ;
        RECT 108.400 91.600 109.200 92.400 ;
        RECT 108.500 90.400 109.100 91.600 ;
        RECT 108.400 89.600 109.200 90.400 ;
        RECT 95.600 81.600 96.400 82.400 ;
        RECT 108.400 82.300 109.200 82.400 ;
        RECT 110.100 82.300 110.700 107.600 ;
        RECT 111.700 98.400 112.300 107.600 ;
        RECT 114.800 104.200 115.600 115.800 ;
        RECT 116.500 114.400 117.100 145.700 ;
        RECT 118.000 126.200 118.800 137.800 ;
        RECT 119.600 135.600 120.400 136.400 ;
        RECT 119.700 118.400 120.300 135.600 ;
        RECT 121.200 130.200 122.000 135.800 ;
        RECT 122.800 135.600 123.600 136.400 ;
        RECT 130.900 134.400 131.500 167.600 ;
        RECT 145.200 166.200 146.000 177.800 ;
        RECT 146.800 173.600 147.600 174.400 ;
        RECT 146.900 172.400 147.500 173.600 ;
        RECT 146.800 171.600 147.600 172.400 ;
        RECT 153.200 171.800 154.000 172.600 ;
        RECT 132.400 151.600 133.200 152.400 ;
        RECT 150.000 151.600 150.800 152.400 ;
        RECT 132.500 146.400 133.100 151.600 ;
        RECT 137.200 149.600 138.000 150.400 ;
        RECT 138.800 149.600 139.600 150.400 ;
        RECT 145.200 149.600 146.000 150.400 ;
        RECT 146.800 149.600 147.600 150.400 ;
        RECT 132.400 145.600 133.200 146.400 ;
        RECT 137.300 144.400 137.900 149.600 ;
        RECT 138.900 148.400 139.500 149.600 ;
        RECT 145.300 148.400 145.900 149.600 ;
        RECT 138.800 147.600 139.600 148.400 ;
        RECT 140.400 147.600 141.200 148.400 ;
        RECT 143.600 147.600 144.400 148.400 ;
        RECT 145.200 147.600 146.000 148.400 ;
        RECT 143.600 145.600 144.400 146.400 ;
        RECT 146.900 146.300 147.500 149.600 ;
        RECT 145.300 145.700 147.500 146.300 ;
        RECT 137.200 143.600 138.000 144.400 ;
        RECT 143.600 143.600 144.400 144.400 ;
        RECT 143.700 136.400 144.300 143.600 ;
        RECT 145.300 136.400 145.900 145.700 ;
        RECT 153.300 144.300 153.900 171.800 ;
        RECT 154.800 166.200 155.600 177.800 ;
        RECT 158.000 170.200 158.800 175.800 ;
        RECT 162.800 173.600 163.600 174.400 ;
        RECT 159.600 171.600 160.400 172.400 ;
        RECT 156.400 153.600 157.200 154.400 ;
        RECT 154.800 149.600 155.600 150.400 ;
        RECT 154.800 147.600 155.600 148.400 ;
        RECT 154.900 146.400 155.500 147.600 ;
        RECT 156.500 146.400 157.100 153.600 ;
        RECT 159.700 152.400 160.300 171.600 ;
        RECT 159.600 151.600 160.400 152.400 ;
        RECT 154.800 145.600 155.600 146.400 ;
        RECT 156.400 145.600 157.200 146.400 ;
        RECT 153.300 143.700 155.500 144.300 ;
        RECT 161.200 144.200 162.000 155.800 ;
        RECT 162.900 150.400 163.500 173.600 ;
        RECT 164.400 170.200 165.200 175.800 ;
        RECT 166.000 173.600 166.800 174.400 ;
        RECT 167.600 166.200 168.400 177.800 ;
        RECT 170.800 171.600 171.600 172.400 ;
        RECT 177.200 166.200 178.000 177.800 ;
        RECT 182.000 177.600 182.800 178.400 ;
        RECT 182.100 174.400 182.700 177.600 ;
        RECT 182.000 173.600 182.800 174.400 ;
        RECT 188.400 173.600 189.200 174.400 ;
        RECT 183.600 171.600 184.400 172.400 ;
        RECT 188.500 172.300 189.100 173.600 ;
        RECT 190.000 172.300 190.800 172.400 ;
        RECT 188.500 171.700 190.800 172.300 ;
        RECT 190.000 171.600 190.800 171.700 ;
        RECT 164.400 151.600 165.200 152.400 ;
        RECT 162.800 149.600 163.600 150.400 ;
        RECT 154.900 138.400 155.500 143.700 ;
        RECT 146.800 137.600 147.600 138.400 ;
        RECT 154.800 137.600 155.600 138.400 ;
        RECT 146.900 136.400 147.500 137.600 ;
        RECT 132.400 135.600 133.200 136.400 ;
        RECT 143.600 135.600 144.400 136.400 ;
        RECT 145.200 135.600 146.000 136.400 ;
        RECT 146.800 135.600 147.600 136.400 ;
        RECT 150.000 135.600 150.800 136.400 ;
        RECT 156.400 135.600 157.200 136.400 ;
        RECT 161.200 135.600 162.000 136.400 ;
        RECT 130.800 133.600 131.600 134.400 ;
        RECT 130.900 132.400 131.500 133.600 ;
        RECT 122.800 131.600 123.600 132.400 ;
        RECT 126.000 131.600 126.800 132.400 ;
        RECT 130.800 131.600 131.600 132.400 ;
        RECT 126.100 128.400 126.700 131.600 ;
        RECT 132.500 130.400 133.100 135.600 ;
        RECT 135.600 133.600 136.400 134.400 ;
        RECT 137.200 133.600 138.000 134.400 ;
        RECT 135.700 132.400 136.300 133.600 ;
        RECT 137.300 132.400 137.900 133.600 ;
        RECT 135.600 131.600 136.400 132.400 ;
        RECT 137.200 131.600 138.000 132.400 ;
        RECT 127.600 129.600 128.400 130.400 ;
        RECT 132.400 129.600 133.200 130.400 ;
        RECT 126.000 127.600 126.800 128.400 ;
        RECT 130.800 127.600 131.600 128.400 ;
        RECT 138.800 127.600 139.600 128.400 ;
        RECT 129.200 123.600 130.000 124.400 ;
        RECT 119.600 117.600 120.400 118.400 ;
        RECT 122.800 117.600 123.600 118.400 ;
        RECT 116.400 113.600 117.200 114.400 ;
        RECT 119.600 113.600 120.400 114.400 ;
        RECT 118.000 106.200 118.800 111.800 ;
        RECT 119.700 110.400 120.300 113.600 ;
        RECT 119.600 109.600 120.400 110.400 ;
        RECT 122.900 106.400 123.500 117.600 ;
        RECT 122.800 105.600 123.600 106.400 ;
        RECT 124.400 106.200 125.200 111.800 ;
        RECT 126.000 109.600 126.800 110.400 ;
        RECT 126.100 108.400 126.700 109.600 ;
        RECT 126.000 107.600 126.800 108.400 ;
        RECT 126.000 105.600 126.800 106.400 ;
        RECT 121.200 103.600 122.000 104.400 ;
        RECT 122.800 103.600 123.600 104.400 ;
        RECT 121.300 102.400 121.900 103.600 ;
        RECT 121.200 101.600 122.000 102.400 ;
        RECT 122.900 98.400 123.500 103.600 ;
        RECT 111.600 97.600 112.400 98.400 ;
        RECT 122.800 97.600 123.600 98.400 ;
        RECT 114.800 95.600 115.600 96.400 ;
        RECT 118.000 95.600 118.800 96.400 ;
        RECT 124.400 96.300 125.200 96.400 ;
        RECT 126.100 96.300 126.700 105.600 ;
        RECT 127.600 104.200 128.400 115.800 ;
        RECT 129.300 114.400 129.900 123.600 ;
        RECT 129.200 113.600 130.000 114.400 ;
        RECT 129.200 111.600 130.000 112.400 ;
        RECT 129.300 110.200 129.900 111.600 ;
        RECT 129.200 109.400 130.000 110.200 ;
        RECT 137.200 104.200 138.000 115.800 ;
        RECT 138.900 114.400 139.500 127.600 ;
        RECT 146.900 118.400 147.500 135.600 ;
        RECT 150.100 132.400 150.700 135.600 ;
        RECT 161.300 134.400 161.900 135.600 ;
        RECT 164.500 134.400 165.100 151.600 ;
        RECT 166.000 149.600 166.800 150.400 ;
        RECT 170.800 144.200 171.600 155.800 ;
        RECT 172.400 149.600 173.200 150.400 ;
        RECT 172.500 142.300 173.100 149.600 ;
        RECT 174.000 146.200 174.800 151.800 ;
        RECT 175.600 146.200 176.400 151.800 ;
        RECT 178.800 144.200 179.600 155.800 ;
        RECT 180.400 149.400 181.200 150.400 ;
        RECT 188.400 144.200 189.200 155.800 ;
        RECT 193.200 143.600 194.000 144.400 ;
        RECT 193.300 142.400 193.900 143.600 ;
        RECT 170.900 141.700 173.100 142.300 ;
        RECT 170.900 138.400 171.500 141.700 ;
        RECT 174.000 141.600 174.800 142.400 ;
        RECT 193.200 141.600 194.000 142.400 ;
        RECT 170.800 137.600 171.600 138.400 ;
        RECT 153.200 133.600 154.000 134.400 ;
        RECT 156.400 133.600 157.200 134.400 ;
        RECT 159.600 133.600 160.400 134.400 ;
        RECT 161.200 133.600 162.000 134.400 ;
        RECT 164.400 133.600 165.200 134.400 ;
        RECT 166.000 133.600 166.800 134.400 ;
        RECT 172.400 133.600 173.200 134.400 ;
        RECT 156.500 132.400 157.100 133.600 ;
        RECT 159.700 132.400 160.300 133.600 ;
        RECT 150.000 131.600 150.800 132.400 ;
        RECT 151.600 131.600 152.400 132.400 ;
        RECT 156.400 131.600 157.200 132.400 ;
        RECT 159.600 131.600 160.400 132.400 ;
        RECT 159.600 129.600 160.400 130.400 ;
        RECT 162.800 130.300 163.600 130.400 ;
        RECT 164.500 130.300 165.100 133.600 ;
        RECT 162.800 129.700 165.100 130.300 ;
        RECT 162.800 129.600 163.600 129.700 ;
        RECT 146.800 117.600 147.600 118.400 ;
        RECT 138.800 113.600 139.600 114.400 ;
        RECT 146.800 111.600 147.600 112.400 ;
        RECT 154.800 111.600 155.600 112.400 ;
        RECT 146.900 108.400 147.500 111.600 ;
        RECT 154.900 108.400 155.500 111.600 ;
        RECT 159.700 110.400 160.300 129.600 ;
        RECT 156.400 109.600 157.200 110.400 ;
        RECT 159.600 109.600 160.400 110.400 ;
        RECT 146.800 107.600 147.600 108.400 ;
        RECT 154.800 107.600 155.600 108.400 ;
        RECT 143.600 105.600 144.400 106.400 ;
        RECT 145.200 103.600 146.000 104.400 ;
        RECT 142.000 101.600 142.800 102.400 ;
        RECT 137.200 97.600 138.000 98.400 ;
        RECT 137.300 96.400 137.900 97.600 ;
        RECT 124.400 95.700 126.700 96.300 ;
        RECT 124.400 95.600 125.200 95.700 ;
        RECT 137.200 95.600 138.000 96.400 ;
        RECT 114.800 93.600 115.600 94.400 ;
        RECT 114.800 87.600 115.600 88.400 ;
        RECT 108.400 81.700 110.700 82.300 ;
        RECT 108.400 81.600 109.200 81.700 ;
        RECT 94.000 71.600 94.800 72.400 ;
        RECT 60.400 69.600 61.200 70.400 ;
        RECT 73.200 69.600 74.000 70.400 ;
        RECT 89.200 69.600 90.000 70.400 ;
        RECT 70.000 63.600 70.800 64.400 ;
        RECT 26.800 53.200 27.600 54.000 ;
        RECT 31.600 53.600 32.400 54.400 ;
        RECT 47.600 53.600 48.400 54.400 ;
        RECT 50.800 50.200 51.600 55.800 ;
        RECT 52.400 53.600 53.200 54.400 ;
        RECT 54.000 46.200 54.800 57.800 ;
        RECT 57.200 51.600 58.000 52.400 ;
        RECT 63.600 46.200 64.400 57.800 ;
        RECT 70.100 54.400 70.700 63.600 ;
        RECT 79.600 56.300 80.400 56.400 ;
        RECT 79.600 55.700 81.900 56.300 ;
        RECT 79.600 55.600 80.400 55.700 ;
        RECT 70.000 53.600 70.800 54.400 ;
        RECT 68.400 43.600 69.200 44.400 ;
        RECT 70.100 36.400 70.700 53.600 ;
        RECT 81.300 52.400 81.900 55.700 ;
        RECT 89.200 55.600 90.000 56.400 ;
        RECT 82.800 53.600 83.600 54.400 ;
        RECT 86.000 53.600 86.800 54.400 ;
        RECT 73.200 51.600 74.000 52.400 ;
        RECT 81.200 51.600 82.000 52.400 ;
        RECT 73.200 49.600 74.000 50.400 ;
        RECT 73.300 38.400 73.900 49.600 ;
        RECT 81.300 44.400 81.900 51.600 ;
        RECT 81.200 43.600 82.000 44.400 ;
        RECT 73.200 37.600 74.000 38.400 ;
        RECT 20.400 35.600 21.200 36.400 ;
        RECT 31.600 35.600 32.400 36.400 ;
        RECT 42.800 35.600 43.600 36.400 ;
        RECT 70.000 35.600 70.800 36.400 ;
        RECT 20.500 32.400 21.100 35.600 ;
        RECT 31.700 32.400 32.300 35.600 ;
        RECT 42.900 32.400 43.500 35.600 ;
        RECT 68.400 33.600 69.200 34.400 ;
        RECT 71.600 33.600 72.400 34.400 ;
        RECT 73.300 32.400 73.900 37.600 ;
        RECT 17.200 27.600 18.000 28.400 ;
        RECT 4.500 12.400 5.100 23.600 ;
        RECT 6.000 17.600 6.800 18.400 ;
        RECT 4.400 11.600 5.200 12.400 ;
        RECT 10.800 6.200 11.600 17.800 ;
        RECT 17.300 14.400 17.900 27.600 ;
        RECT 18.800 26.200 19.600 31.800 ;
        RECT 20.400 31.600 21.200 32.400 ;
        RECT 31.600 31.600 32.400 32.400 ;
        RECT 42.800 31.600 43.600 32.400 ;
        RECT 44.400 31.600 45.200 32.400 ;
        RECT 58.800 31.600 59.600 32.400 ;
        RECT 65.200 31.600 66.000 32.400 ;
        RECT 71.600 31.600 72.400 32.400 ;
        RECT 73.200 31.600 74.000 32.400 ;
        RECT 23.600 29.600 24.400 30.400 ;
        RECT 25.200 29.600 26.000 30.400 ;
        RECT 23.700 28.400 24.300 29.600 ;
        RECT 23.600 27.600 24.400 28.400 ;
        RECT 25.200 27.600 26.000 28.400 ;
        RECT 26.800 27.600 27.600 28.400 ;
        RECT 36.400 27.600 37.200 28.400 ;
        RECT 41.200 27.600 42.000 28.400 ;
        RECT 25.300 26.400 25.900 27.600 ;
        RECT 26.900 26.400 27.500 27.600 ;
        RECT 25.200 25.600 26.000 26.400 ;
        RECT 26.800 25.600 27.600 26.400 ;
        RECT 30.000 25.600 30.800 26.400 ;
        RECT 20.400 23.600 21.200 24.400 ;
        RECT 20.500 20.400 21.100 23.600 ;
        RECT 20.400 19.600 21.200 20.400 ;
        RECT 25.200 19.600 26.000 20.400 ;
        RECT 17.200 13.600 18.000 14.400 ;
        RECT 18.800 11.600 19.600 12.600 ;
        RECT 20.400 6.200 21.200 17.800 ;
        RECT 25.300 16.400 25.900 19.600 ;
        RECT 23.600 10.200 24.400 15.800 ;
        RECT 25.200 15.600 26.000 16.400 ;
        RECT 25.200 11.600 26.000 12.400 ;
        RECT 26.900 12.300 27.500 25.600 ;
        RECT 30.100 18.400 30.700 25.600 ;
        RECT 36.500 24.400 37.100 27.600 ;
        RECT 38.000 25.600 38.800 26.400 ;
        RECT 36.400 23.600 37.200 24.400 ;
        RECT 30.000 17.600 30.800 18.400 ;
        RECT 30.100 16.400 30.700 17.600 ;
        RECT 30.000 15.600 30.800 16.400 ;
        RECT 28.400 13.600 29.200 14.400 ;
        RECT 28.500 12.400 29.100 13.600 ;
        RECT 30.100 12.400 30.700 15.600 ;
        RECT 36.500 14.400 37.100 23.600 ;
        RECT 36.400 13.600 37.200 14.400 ;
        RECT 38.100 12.400 38.700 25.600 ;
        RECT 42.800 23.600 43.600 24.400 ;
        RECT 42.900 18.400 43.500 23.600 ;
        RECT 42.800 17.600 43.600 18.400 ;
        RECT 44.500 16.400 45.100 31.600 ;
        RECT 65.300 30.400 65.900 31.600 ;
        RECT 46.000 29.600 46.800 30.400 ;
        RECT 52.400 29.600 53.200 30.400 ;
        RECT 65.200 29.600 66.000 30.400 ;
        RECT 47.600 27.600 48.400 28.400 ;
        RECT 58.800 27.600 59.600 28.400 ;
        RECT 63.600 27.600 64.400 28.400 ;
        RECT 47.600 17.600 48.400 18.400 ;
        RECT 47.700 16.400 48.300 17.600 ;
        RECT 39.600 15.600 40.400 16.400 ;
        RECT 44.400 15.600 45.200 16.400 ;
        RECT 47.600 15.600 48.400 16.400 ;
        RECT 39.700 14.400 40.300 15.600 ;
        RECT 39.600 13.600 40.400 14.400 ;
        RECT 28.400 12.300 29.200 12.400 ;
        RECT 26.900 11.700 29.200 12.300 ;
        RECT 28.400 11.600 29.200 11.700 ;
        RECT 30.000 11.600 30.800 12.400 ;
        RECT 31.600 11.600 32.400 12.400 ;
        RECT 38.000 11.600 38.800 12.400 ;
        RECT 52.400 11.600 53.200 12.400 ;
        RECT 54.000 10.200 54.800 15.800 ;
        RECT 55.600 13.600 56.400 14.400 ;
        RECT 57.200 6.200 58.000 17.800 ;
        RECT 63.700 16.400 64.300 27.600 ;
        RECT 71.700 18.400 72.300 31.600 ;
        RECT 73.200 29.600 74.000 30.400 ;
        RECT 79.600 29.600 80.400 30.400 ;
        RECT 73.300 26.400 73.900 29.600 ;
        RECT 81.300 28.400 81.900 43.600 ;
        RECT 82.900 30.400 83.500 53.600 ;
        RECT 86.100 52.400 86.700 53.600 ;
        RECT 84.400 51.600 85.200 52.400 ;
        RECT 86.000 51.600 86.800 52.400 ;
        RECT 84.500 48.400 85.100 51.600 ;
        RECT 94.100 50.400 94.700 71.600 ;
        RECT 97.200 69.600 98.000 70.400 ;
        RECT 98.800 69.600 99.600 70.400 ;
        RECT 105.200 69.600 106.000 70.400 ;
        RECT 95.600 67.600 96.400 68.400 ;
        RECT 95.700 66.400 96.300 67.600 ;
        RECT 95.600 65.600 96.400 66.400 ;
        RECT 97.300 64.400 97.900 69.600 ;
        RECT 98.900 68.400 99.500 69.600 ;
        RECT 98.800 67.600 99.600 68.400 ;
        RECT 102.000 67.600 102.800 68.400 ;
        RECT 105.200 67.600 106.000 68.400 ;
        RECT 100.400 65.600 101.200 66.400 ;
        RECT 105.300 64.400 105.900 67.600 ;
        RECT 106.800 66.200 107.600 71.800 ;
        RECT 108.500 68.400 109.100 81.600 ;
        RECT 108.400 67.600 109.200 68.400 ;
        RECT 97.200 63.600 98.000 64.400 ;
        RECT 105.200 63.600 106.000 64.400 ;
        RECT 110.000 64.200 110.800 75.800 ;
        RECT 111.600 69.400 112.400 70.200 ;
        RECT 111.700 68.400 112.300 69.400 ;
        RECT 111.600 67.600 112.400 68.400 ;
        RECT 105.300 58.400 105.900 63.600 ;
        RECT 105.200 57.600 106.000 58.400 ;
        RECT 110.000 55.600 110.800 56.400 ;
        RECT 89.200 49.600 90.000 50.400 ;
        RECT 94.000 49.600 94.800 50.400 ;
        RECT 105.200 49.600 106.000 50.400 ;
        RECT 84.400 47.600 85.200 48.400 ;
        RECT 82.800 29.600 83.600 30.400 ;
        RECT 84.500 28.400 85.100 47.600 ;
        RECT 89.300 30.400 89.900 49.600 ;
        RECT 94.100 32.400 94.700 49.600 ;
        RECT 105.300 48.400 105.900 49.600 ;
        RECT 105.200 47.600 106.000 48.400 ;
        RECT 102.000 43.600 102.800 44.400 ;
        RECT 102.100 32.400 102.700 43.600 ;
        RECT 94.000 31.600 94.800 32.400 ;
        RECT 98.800 31.600 99.600 32.400 ;
        RECT 102.000 31.600 102.800 32.400 ;
        RECT 114.900 32.300 115.500 87.600 ;
        RECT 116.400 53.600 117.200 54.400 ;
        RECT 116.400 51.600 117.200 52.400 ;
        RECT 116.500 44.300 117.100 51.600 ;
        RECT 118.100 46.400 118.700 95.600 ;
        RECT 121.200 93.600 122.000 94.400 ;
        RECT 129.200 93.600 130.000 94.400 ;
        RECT 134.000 93.600 134.800 94.400 ;
        RECT 129.300 92.400 129.900 93.600 ;
        RECT 137.300 92.400 137.900 95.600 ;
        RECT 142.100 94.400 142.700 101.600 ;
        RECT 143.600 99.600 144.400 100.400 ;
        RECT 143.700 96.400 144.300 99.600 ;
        RECT 145.300 96.400 145.900 103.600 ;
        RECT 143.600 95.600 144.400 96.400 ;
        RECT 145.200 95.600 146.000 96.400 ;
        RECT 143.700 94.400 144.300 95.600 ;
        RECT 142.000 93.600 142.800 94.400 ;
        RECT 143.600 93.600 144.400 94.400 ;
        RECT 145.200 93.600 146.000 94.400 ;
        RECT 119.600 91.600 120.400 92.400 ;
        RECT 126.000 91.600 126.800 92.400 ;
        RECT 129.200 91.600 130.000 92.400 ;
        RECT 130.800 91.600 131.600 92.400 ;
        RECT 132.400 91.600 133.200 92.400 ;
        RECT 137.200 91.600 138.000 92.400 ;
        RECT 127.600 87.600 128.400 88.400 ;
        RECT 127.700 80.400 128.300 87.600 ;
        RECT 132.500 80.400 133.100 91.600 ;
        RECT 146.900 90.400 147.500 107.600 ;
        RECT 148.400 95.600 149.200 96.400 ;
        RECT 153.200 95.600 154.000 96.400 ;
        RECT 148.500 94.400 149.100 95.600 ;
        RECT 156.500 94.400 157.100 109.600 ;
        RECT 162.900 108.400 163.500 129.600 ;
        RECT 166.100 118.400 166.700 133.600 ;
        RECT 174.100 132.400 174.700 141.600 ;
        RECT 174.000 131.600 174.800 132.400 ;
        RECT 167.600 129.600 168.400 130.400 ;
        RECT 166.000 117.600 166.800 118.400 ;
        RECT 170.800 115.600 171.600 116.400 ;
        RECT 170.900 112.400 171.500 115.600 ;
        RECT 172.400 113.600 173.200 114.400 ;
        RECT 167.600 111.600 168.400 112.400 ;
        RECT 169.200 111.600 170.000 112.400 ;
        RECT 170.800 111.600 171.600 112.400 ;
        RECT 164.400 109.600 165.200 110.400 ;
        RECT 162.800 107.600 163.600 108.400 ;
        RECT 164.400 107.600 165.200 108.400 ;
        RECT 164.500 106.400 165.100 107.600 ;
        RECT 167.700 106.400 168.300 111.600 ;
        RECT 164.400 105.600 165.200 106.400 ;
        RECT 167.600 105.600 168.400 106.400 ;
        RECT 169.300 98.400 169.900 111.600 ;
        RECT 170.800 109.600 171.600 110.400 ;
        RECT 170.900 100.400 171.500 109.600 ;
        RECT 172.500 104.400 173.100 113.600 ;
        RECT 174.100 108.400 174.700 131.600 ;
        RECT 175.600 130.200 176.400 135.800 ;
        RECT 177.200 133.600 178.000 134.400 ;
        RECT 177.300 128.400 177.900 133.600 ;
        RECT 177.200 127.600 178.000 128.400 ;
        RECT 178.800 126.200 179.600 137.800 ;
        RECT 183.600 131.600 184.400 132.400 ;
        RECT 183.700 124.300 184.300 131.600 ;
        RECT 188.400 126.200 189.200 137.800 ;
        RECT 183.700 123.700 185.900 124.300 ;
        RECT 185.300 118.400 185.900 123.700 ;
        RECT 193.200 123.600 194.000 124.400 ;
        RECT 185.200 117.600 186.000 118.400 ;
        RECT 180.400 109.600 181.200 110.400 ;
        RECT 188.400 109.600 189.200 110.400 ;
        RECT 174.000 107.600 174.800 108.400 ;
        RECT 175.600 107.600 176.400 108.400 ;
        RECT 175.700 106.300 176.300 107.600 ;
        RECT 174.100 105.700 176.300 106.300 ;
        RECT 172.400 103.600 173.200 104.400 ;
        RECT 170.800 99.600 171.600 100.400 ;
        RECT 159.600 97.600 160.400 98.400 ;
        RECT 169.200 97.600 170.000 98.400 ;
        RECT 159.700 96.400 160.300 97.600 ;
        RECT 159.600 95.600 160.400 96.400 ;
        RECT 148.400 93.600 149.200 94.400 ;
        RECT 151.600 93.600 152.400 94.400 ;
        RECT 156.400 93.600 157.200 94.400 ;
        RECT 158.000 93.600 158.800 94.400 ;
        RECT 166.000 93.600 166.800 94.400 ;
        RECT 156.500 92.400 157.100 93.600 ;
        RECT 158.100 92.400 158.700 93.600 ;
        RECT 172.500 92.400 173.100 103.600 ;
        RECT 174.100 98.400 174.700 105.700 ;
        RECT 180.500 102.400 181.100 109.600 ;
        RECT 188.500 108.400 189.100 109.600 ;
        RECT 188.400 107.600 189.200 108.400 ;
        RECT 193.300 106.400 193.900 123.600 ;
        RECT 188.400 105.600 189.200 106.400 ;
        RECT 193.200 105.600 194.000 106.400 ;
        RECT 180.400 101.600 181.200 102.400 ;
        RECT 183.600 99.600 184.400 100.400 ;
        RECT 174.000 97.600 174.800 98.400 ;
        RECT 182.000 95.600 182.800 96.400 ;
        RECT 150.000 91.600 150.800 92.400 ;
        RECT 156.400 91.600 157.200 92.400 ;
        RECT 158.000 91.600 158.800 92.400 ;
        RECT 164.400 91.600 165.200 92.400 ;
        RECT 172.400 91.600 173.200 92.400 ;
        RECT 146.800 89.600 147.600 90.400 ;
        RECT 153.200 83.600 154.000 84.400 ;
        RECT 122.800 79.600 123.600 80.400 ;
        RECT 127.600 79.600 128.400 80.400 ;
        RECT 132.400 79.600 133.200 80.400 ;
        RECT 119.600 64.200 120.400 75.800 ;
        RECT 122.900 58.400 123.500 79.600 ;
        RECT 153.300 74.400 153.900 83.600 ;
        RECT 126.000 73.600 126.800 74.400 ;
        RECT 153.200 73.600 154.000 74.400 ;
        RECT 126.100 66.400 126.700 73.600 ;
        RECT 134.000 71.600 134.800 72.400 ;
        RECT 146.800 71.600 147.600 72.400 ;
        RECT 153.200 72.300 154.000 72.400 ;
        RECT 151.700 71.700 154.000 72.300 ;
        RECT 127.600 69.600 128.400 70.400 ;
        RECT 130.800 69.600 131.600 70.400 ;
        RECT 138.800 69.600 139.600 70.400 ;
        RECT 142.000 69.600 142.800 70.400 ;
        RECT 145.200 69.600 146.000 70.400 ;
        RECT 126.000 65.600 126.800 66.400 ;
        RECT 130.900 64.400 131.500 69.600 ;
        RECT 140.400 68.300 141.200 68.400 ;
        RECT 140.400 67.700 142.700 68.300 ;
        RECT 140.400 67.600 141.200 67.700 ;
        RECT 129.200 63.600 130.000 64.400 ;
        RECT 130.800 63.600 131.600 64.400 ;
        RECT 122.800 57.600 123.600 58.400 ;
        RECT 127.600 57.600 128.400 58.400 ;
        RECT 122.800 55.600 123.600 56.400 ;
        RECT 122.900 52.400 123.500 55.600 ;
        RECT 127.700 54.400 128.300 57.600 ;
        RECT 127.600 53.600 128.400 54.400 ;
        RECT 129.300 52.400 129.900 63.600 ;
        RECT 138.800 57.600 139.600 58.400 ;
        RECT 138.900 56.400 139.500 57.600 ;
        RECT 142.100 56.400 142.700 67.700 ;
        RECT 150.000 67.600 150.800 68.400 ;
        RECT 150.100 64.400 150.700 67.600 ;
        RECT 151.700 66.400 152.300 71.700 ;
        RECT 153.200 71.600 154.000 71.700 ;
        RECT 151.600 65.600 152.400 66.400 ;
        RECT 150.000 63.600 150.800 64.400 ;
        RECT 145.200 57.600 146.000 58.400 ;
        RECT 146.800 57.600 147.600 58.400 ;
        RECT 138.800 55.600 139.600 56.400 ;
        RECT 142.000 55.600 142.800 56.400 ;
        RECT 143.600 55.600 144.400 56.400 ;
        RECT 143.700 54.400 144.300 55.600 ;
        RECT 143.600 53.600 144.400 54.400 ;
        RECT 121.200 51.600 122.000 52.400 ;
        RECT 122.800 51.600 123.600 52.400 ;
        RECT 129.200 51.600 130.000 52.400 ;
        RECT 142.000 51.600 142.800 52.400 ;
        RECT 118.000 45.600 118.800 46.400 ;
        RECT 116.500 43.700 118.700 44.300 ;
        RECT 116.400 32.300 117.200 32.400 ;
        RECT 114.900 31.700 117.200 32.300 ;
        RECT 116.400 31.600 117.200 31.700 ;
        RECT 98.900 30.400 99.500 31.600 ;
        RECT 89.200 29.600 90.000 30.400 ;
        RECT 90.800 29.600 91.600 30.400 ;
        RECT 98.800 29.600 99.600 30.400 ;
        RECT 102.000 29.600 102.800 30.400 ;
        RECT 108.400 29.600 109.200 30.400 ;
        RECT 113.200 29.600 114.000 30.400 ;
        RECT 89.300 28.400 89.900 29.600 ;
        RECT 90.900 28.400 91.500 29.600 ;
        RECT 98.900 28.400 99.500 29.600 ;
        RECT 113.300 28.400 113.900 29.600 ;
        RECT 118.100 28.400 118.700 43.700 ;
        RECT 119.600 30.300 120.400 30.400 ;
        RECT 121.300 30.300 121.900 51.600 ;
        RECT 142.100 50.400 142.700 51.600 ;
        RECT 132.400 49.600 133.200 50.400 ;
        RECT 142.000 49.600 142.800 50.400 ;
        RECT 145.200 50.300 146.000 50.400 ;
        RECT 146.900 50.300 147.500 57.600 ;
        RECT 150.100 54.400 150.700 63.600 ;
        RECT 148.400 53.600 149.200 54.400 ;
        RECT 150.000 53.600 150.800 54.400 ;
        RECT 148.500 50.400 149.100 53.600 ;
        RECT 145.200 49.700 147.500 50.300 ;
        RECT 145.200 49.600 146.000 49.700 ;
        RECT 148.400 49.600 149.200 50.400 ;
        RECT 129.200 43.600 130.000 44.400 ;
        RECT 122.800 31.600 123.600 32.400 ;
        RECT 119.600 29.700 121.900 30.300 ;
        RECT 119.600 29.600 120.400 29.700 ;
        RECT 122.900 28.400 123.500 31.600 ;
        RECT 81.200 27.600 82.000 28.400 ;
        RECT 84.400 27.600 85.200 28.400 ;
        RECT 89.200 27.600 90.000 28.400 ;
        RECT 90.800 27.600 91.600 28.400 ;
        RECT 92.400 27.600 93.200 28.400 ;
        RECT 97.200 27.600 98.000 28.400 ;
        RECT 98.800 27.600 99.600 28.400 ;
        RECT 103.600 27.600 104.400 28.400 ;
        RECT 113.200 27.600 114.000 28.400 ;
        RECT 116.400 27.600 117.200 28.400 ;
        RECT 118.000 27.600 118.800 28.400 ;
        RECT 122.800 27.600 123.600 28.400 ;
        RECT 73.200 25.600 74.000 26.400 ;
        RECT 63.600 15.600 64.400 16.400 ;
        RECT 58.800 11.600 59.600 12.600 ;
        RECT 63.700 12.400 64.300 15.600 ;
        RECT 63.600 11.600 64.400 12.400 ;
        RECT 66.800 6.200 67.600 17.800 ;
        RECT 71.600 17.600 72.400 18.400 ;
        RECT 71.700 14.400 72.300 17.600 ;
        RECT 71.600 13.600 72.400 14.400 ;
        RECT 78.000 13.600 78.800 14.400 ;
        RECT 78.100 12.400 78.700 13.600 ;
        RECT 81.300 12.400 81.900 27.600 ;
        RECT 87.600 25.600 88.400 26.400 ;
        RECT 86.000 23.600 86.800 24.400 ;
        RECT 86.100 14.400 86.700 23.600 ;
        RECT 89.300 18.400 89.900 27.600 ;
        RECT 92.500 26.400 93.100 27.600 ;
        RECT 97.300 26.400 97.900 27.600 ;
        RECT 92.400 25.600 93.200 26.400 ;
        RECT 97.200 25.600 98.000 26.400 ;
        RECT 106.800 25.600 107.600 26.400 ;
        RECT 110.000 25.600 110.800 26.400 ;
        RECT 105.200 23.600 106.000 24.400 ;
        RECT 89.200 17.600 90.000 18.400 ;
        RECT 92.400 17.600 93.200 18.400 ;
        RECT 97.200 17.600 98.000 18.400 ;
        RECT 82.800 13.600 83.600 14.400 ;
        RECT 86.000 13.600 86.800 14.400 ;
        RECT 82.900 12.400 83.500 13.600 ;
        RECT 92.500 12.400 93.100 17.600 ;
        RECT 76.400 11.600 77.200 12.400 ;
        RECT 78.000 11.600 78.800 12.400 ;
        RECT 81.200 11.600 82.000 12.400 ;
        RECT 82.800 11.600 83.600 12.400 ;
        RECT 87.600 11.600 88.400 12.400 ;
        RECT 92.400 11.600 93.200 12.400 ;
        RECT 102.000 6.200 102.800 17.800 ;
        RECT 105.300 10.400 105.900 23.600 ;
        RECT 106.800 15.600 107.600 16.400 ;
        RECT 106.900 14.400 107.500 15.600 ;
        RECT 106.800 13.600 107.600 14.400 ;
        RECT 108.400 13.600 109.200 14.400 ;
        RECT 108.500 12.400 109.100 13.600 ;
        RECT 110.100 12.400 110.700 25.600 ;
        RECT 118.100 18.400 118.700 27.600 ;
        RECT 129.300 26.400 129.900 43.600 ;
        RECT 132.400 29.600 133.200 30.400 ;
        RECT 129.200 25.600 130.000 26.400 ;
        RECT 134.000 26.200 134.800 31.800 ;
        RECT 137.200 24.200 138.000 35.800 ;
        RECT 138.800 29.400 139.600 30.400 ;
        RECT 142.000 29.600 142.800 30.400 ;
        RECT 142.100 28.400 142.700 29.600 ;
        RECT 142.000 27.600 142.800 28.400 ;
        RECT 108.400 11.600 109.200 12.400 ;
        RECT 110.000 11.600 110.800 12.400 ;
        RECT 105.200 9.600 106.000 10.400 ;
        RECT 111.600 6.200 112.400 17.800 ;
        RECT 116.400 17.600 117.200 18.400 ;
        RECT 118.000 17.600 118.800 18.400 ;
        RECT 114.800 10.200 115.600 15.800 ;
        RECT 116.500 12.400 117.100 17.600 ;
        RECT 119.600 13.600 120.400 14.400 ;
        RECT 119.700 12.400 120.300 13.600 ;
        RECT 116.400 11.600 117.200 12.400 ;
        RECT 119.600 11.600 120.400 12.400 ;
        RECT 116.500 10.400 117.100 11.600 ;
        RECT 116.400 9.600 117.200 10.400 ;
        RECT 121.200 10.200 122.000 15.800 ;
        RECT 122.800 15.600 123.600 16.400 ;
        RECT 122.900 14.400 123.500 15.600 ;
        RECT 122.800 13.600 123.600 14.400 ;
        RECT 124.400 6.200 125.200 17.800 ;
        RECT 126.000 11.800 126.800 12.600 ;
        RECT 126.100 10.400 126.700 11.800 ;
        RECT 126.000 9.600 126.800 10.400 ;
        RECT 134.000 6.200 134.800 17.800 ;
        RECT 138.800 17.600 139.600 18.400 ;
        RECT 142.100 16.400 142.700 27.600 ;
        RECT 146.800 24.200 147.600 35.800 ;
        RECT 142.000 15.600 142.800 16.400 ;
        RECT 150.100 14.400 150.700 53.600 ;
        RECT 151.700 52.400 152.300 65.600 ;
        RECT 153.200 63.600 154.000 64.400 ;
        RECT 154.800 63.600 155.600 64.400 ;
        RECT 159.600 64.200 160.400 75.800 ;
        RECT 153.300 60.400 153.900 63.600 ;
        RECT 159.600 61.600 160.400 62.400 ;
        RECT 153.200 59.600 154.000 60.400 ;
        RECT 158.000 55.600 158.800 56.400 ;
        RECT 158.000 53.600 158.800 54.400 ;
        RECT 158.100 52.400 158.700 53.600 ;
        RECT 151.600 51.600 152.400 52.400 ;
        RECT 153.200 51.600 154.000 52.400 ;
        RECT 158.000 51.600 158.800 52.400 ;
        RECT 151.700 28.400 152.300 51.600 ;
        RECT 153.300 38.400 153.900 51.600 ;
        RECT 154.800 49.600 155.600 50.400 ;
        RECT 158.000 47.600 158.800 48.400 ;
        RECT 153.200 37.600 154.000 38.400 ;
        RECT 151.600 27.600 152.400 28.400 ;
        RECT 154.800 27.600 155.600 28.400 ;
        RECT 151.600 23.600 152.400 24.400 ;
        RECT 150.000 13.600 150.800 14.400 ;
        RECT 150.000 12.300 150.800 12.400 ;
        RECT 151.700 12.300 152.300 23.600 ;
        RECT 154.900 12.400 155.500 27.600 ;
        RECT 158.000 24.200 158.800 35.800 ;
        RECT 159.700 30.400 160.300 61.600 ;
        RECT 164.500 58.400 165.100 91.600 ;
        RECT 182.100 90.300 182.700 95.600 ;
        RECT 183.700 92.400 184.300 99.600 ;
        RECT 188.500 98.400 189.100 105.600 ;
        RECT 191.600 99.600 192.400 100.400 ;
        RECT 188.400 97.600 189.200 98.400 ;
        RECT 188.500 92.400 189.100 97.600 ;
        RECT 183.600 91.600 184.400 92.400 ;
        RECT 188.400 91.600 189.200 92.400 ;
        RECT 182.100 89.700 184.300 90.300 ;
        RECT 180.400 83.600 181.200 84.400 ;
        RECT 166.000 69.600 166.800 70.400 ;
        RECT 167.600 65.600 168.400 66.400 ;
        RECT 167.700 62.400 168.300 65.600 ;
        RECT 169.200 64.200 170.000 75.800 ;
        RECT 172.400 66.200 173.200 71.800 ;
        RECT 174.000 66.200 174.800 71.800 ;
        RECT 175.600 67.600 176.400 68.400 ;
        RECT 175.700 62.400 176.300 67.600 ;
        RECT 177.200 64.200 178.000 75.800 ;
        RECT 178.800 73.600 179.600 74.400 ;
        RECT 178.900 70.200 179.500 73.600 ;
        RECT 178.800 69.400 179.600 70.200 ;
        RECT 167.600 61.600 168.400 62.400 ;
        RECT 175.600 61.600 176.400 62.400 ;
        RECT 169.200 59.600 170.000 60.400 ;
        RECT 164.400 57.600 165.200 58.400 ;
        RECT 169.300 56.400 169.900 59.600 ;
        RECT 174.000 57.600 174.800 58.400 ;
        RECT 180.500 58.300 181.100 83.600 ;
        RECT 180.500 57.700 182.700 58.300 ;
        RECT 169.200 55.600 170.000 56.400 ;
        RECT 172.400 55.600 173.200 56.400 ;
        RECT 180.400 55.600 181.200 56.400 ;
        RECT 166.000 53.600 166.800 54.400 ;
        RECT 166.100 52.400 166.700 53.600 ;
        RECT 172.500 52.400 173.100 55.600 ;
        RECT 180.400 53.600 181.200 54.400 ;
        RECT 166.000 51.600 166.800 52.400 ;
        RECT 169.200 51.600 170.000 52.400 ;
        RECT 172.400 51.600 173.200 52.400 ;
        RECT 177.200 51.600 178.000 52.400 ;
        RECT 178.800 51.600 179.600 52.400 ;
        RECT 167.600 50.300 168.400 50.400 ;
        RECT 169.300 50.300 169.900 51.600 ;
        RECT 167.600 49.700 169.900 50.300 ;
        RECT 177.300 50.300 177.900 51.600 ;
        RECT 178.900 50.400 179.500 51.600 ;
        RECT 178.800 50.300 179.600 50.400 ;
        RECT 177.300 49.700 179.600 50.300 ;
        RECT 167.600 49.600 168.400 49.700 ;
        RECT 178.800 49.600 179.600 49.700 ;
        RECT 164.400 47.600 165.200 48.400 ;
        RECT 161.200 43.600 162.000 44.400 ;
        RECT 159.600 29.600 160.400 30.400 ;
        RECT 159.600 25.600 160.400 26.400 ;
        RECT 159.700 16.400 160.300 25.600 ;
        RECT 159.600 15.600 160.400 16.400 ;
        RECT 159.600 13.600 160.400 14.400 ;
        RECT 159.700 12.400 160.300 13.600 ;
        RECT 161.300 12.400 161.900 43.600 ;
        RECT 166.000 29.400 166.800 30.400 ;
        RECT 167.600 24.200 168.400 35.800 ;
        RECT 170.800 26.200 171.600 31.800 ;
        RECT 172.400 26.200 173.200 31.800 ;
        RECT 175.600 24.200 176.400 35.800 ;
        RECT 178.800 29.600 179.600 30.400 ;
        RECT 180.400 29.600 181.200 30.400 ;
        RECT 178.900 28.400 179.500 29.600 ;
        RECT 178.800 27.600 179.600 28.400 ;
        RECT 180.500 18.400 181.100 29.600 ;
        RECT 180.400 17.600 181.200 18.400 ;
        RECT 182.100 16.400 182.700 57.700 ;
        RECT 183.700 54.400 184.300 89.700 ;
        RECT 191.700 78.400 192.300 99.600 ;
        RECT 191.600 77.600 192.400 78.400 ;
        RECT 186.800 64.200 187.600 75.800 ;
        RECT 183.600 53.600 184.400 54.400 ;
        RECT 183.700 38.400 184.300 53.600 ;
        RECT 190.000 51.600 190.800 52.400 ;
        RECT 183.600 37.600 184.400 38.400 ;
        RECT 190.000 37.600 190.800 38.400 ;
        RECT 185.200 24.200 186.000 35.800 ;
        RECT 188.400 27.600 189.200 28.400 ;
        RECT 186.800 25.600 187.600 26.400 ;
        RECT 186.900 16.400 187.500 25.600 ;
        RECT 188.500 18.400 189.100 27.600 ;
        RECT 188.400 17.600 189.200 18.400 ;
        RECT 164.400 15.600 165.200 16.400 ;
        RECT 167.600 15.600 168.400 16.400 ;
        RECT 174.000 15.600 174.800 16.400 ;
        RECT 182.000 15.600 182.800 16.400 ;
        RECT 186.800 15.600 187.600 16.400 ;
        RECT 190.000 15.600 190.800 16.400 ;
        RECT 167.700 12.400 168.300 15.600 ;
        RECT 190.100 14.400 190.700 15.600 ;
        RECT 169.200 13.600 170.000 14.400 ;
        RECT 175.600 13.600 176.400 14.400 ;
        RECT 178.800 13.600 179.600 14.400 ;
        RECT 185.200 13.600 186.000 14.400 ;
        RECT 190.000 13.600 190.800 14.400 ;
        RECT 191.600 13.600 192.400 14.400 ;
        RECT 191.700 12.400 192.300 13.600 ;
        RECT 150.000 11.700 152.300 12.300 ;
        RECT 150.000 11.600 150.800 11.700 ;
        RECT 154.800 11.600 155.600 12.400 ;
        RECT 159.600 11.600 160.400 12.400 ;
        RECT 161.200 11.600 162.000 12.400 ;
        RECT 167.600 11.600 168.400 12.400 ;
        RECT 172.400 11.600 173.200 12.400 ;
        RECT 183.600 11.600 184.400 12.400 ;
        RECT 191.600 11.600 192.400 12.400 ;
      LAYER via2 ;
        RECT 33.200 149.600 34.000 150.400 ;
        RECT 14.000 29.600 14.800 30.400 ;
        RECT 180.400 149.600 181.200 150.400 ;
        RECT 138.800 29.600 139.600 30.400 ;
        RECT 166.000 29.600 166.800 30.400 ;
      LAYER metal3 ;
        RECT 26.800 174.300 27.600 174.400 ;
        RECT 41.200 174.300 42.000 174.400 ;
        RECT 26.800 173.700 42.000 174.300 ;
        RECT 26.800 173.600 27.600 173.700 ;
        RECT 41.200 173.600 42.000 173.700 ;
        RECT 94.000 174.300 94.800 174.400 ;
        RECT 113.200 174.300 114.000 174.400 ;
        RECT 146.800 174.300 147.600 174.400 ;
        RECT 162.800 174.300 163.600 174.400 ;
        RECT 166.000 174.300 166.800 174.400 ;
        RECT 94.000 173.700 166.800 174.300 ;
        RECT 94.000 173.600 94.800 173.700 ;
        RECT 113.200 173.600 114.000 173.700 ;
        RECT 146.800 173.600 147.600 173.700 ;
        RECT 162.800 173.600 163.600 173.700 ;
        RECT 166.000 173.600 166.800 173.700 ;
        RECT 182.000 174.300 182.800 174.400 ;
        RECT 188.400 174.300 189.200 174.400 ;
        RECT 182.000 173.700 189.200 174.300 ;
        RECT 182.000 173.600 182.800 173.700 ;
        RECT 188.400 173.600 189.200 173.700 ;
        RECT 97.200 172.300 98.000 172.400 ;
        RECT 100.400 172.300 101.200 172.400 ;
        RECT 97.200 171.700 101.200 172.300 ;
        RECT 97.200 171.600 98.000 171.700 ;
        RECT 100.400 171.600 101.200 171.700 ;
        RECT 170.800 172.300 171.600 172.400 ;
        RECT 183.600 172.300 184.400 172.400 ;
        RECT 170.800 171.700 184.400 172.300 ;
        RECT 170.800 171.600 171.600 171.700 ;
        RECT 183.600 171.600 184.400 171.700 ;
        RECT 90.800 170.300 91.600 170.400 ;
        RECT 100.400 170.300 101.200 170.400 ;
        RECT 90.800 169.700 101.200 170.300 ;
        RECT 90.800 169.600 91.600 169.700 ;
        RECT 100.400 169.600 101.200 169.700 ;
        RECT 130.800 168.300 131.600 168.400 ;
        RECT 140.400 168.300 141.200 168.400 ;
        RECT 130.800 167.700 141.200 168.300 ;
        RECT 130.800 167.600 131.600 167.700 ;
        RECT 140.400 167.600 141.200 167.700 ;
        RECT 28.400 166.300 29.200 166.400 ;
        RECT 39.600 166.300 40.400 166.400 ;
        RECT 28.400 165.700 40.400 166.300 ;
        RECT 28.400 165.600 29.200 165.700 ;
        RECT 39.600 165.600 40.400 165.700 ;
        RECT 46.000 166.300 46.800 166.400 ;
        RECT 70.000 166.300 70.800 166.400 ;
        RECT 46.000 165.700 70.800 166.300 ;
        RECT 46.000 165.600 46.800 165.700 ;
        RECT 70.000 165.600 70.800 165.700 ;
        RECT 73.200 166.300 74.000 166.400 ;
        RECT 78.000 166.300 78.800 166.400 ;
        RECT 73.200 165.700 78.800 166.300 ;
        RECT 73.200 165.600 74.000 165.700 ;
        RECT 78.000 165.600 78.800 165.700 ;
        RECT 15.600 160.300 16.400 160.400 ;
        RECT 23.600 160.300 24.400 160.400 ;
        RECT 34.800 160.300 35.600 160.400 ;
        RECT 15.600 159.700 35.600 160.300 ;
        RECT 15.600 159.600 16.400 159.700 ;
        RECT 23.600 159.600 24.400 159.700 ;
        RECT 34.800 159.600 35.600 159.700 ;
        RECT 126.000 160.300 126.800 160.400 ;
        RECT 129.200 160.300 130.000 160.400 ;
        RECT 126.000 159.700 130.000 160.300 ;
        RECT 126.000 159.600 126.800 159.700 ;
        RECT 129.200 159.600 130.000 159.700 ;
        RECT 58.800 152.300 59.600 152.400 ;
        RECT 65.200 152.300 66.000 152.400 ;
        RECT 68.400 152.300 69.200 152.400 ;
        RECT 74.800 152.300 75.600 152.400 ;
        RECT 58.800 151.700 75.600 152.300 ;
        RECT 58.800 151.600 59.600 151.700 ;
        RECT 65.200 151.600 66.000 151.700 ;
        RECT 68.400 151.600 69.200 151.700 ;
        RECT 74.800 151.600 75.600 151.700 ;
        RECT 122.800 152.300 123.600 152.400 ;
        RECT 150.000 152.300 150.800 152.400 ;
        RECT 164.400 152.300 165.200 152.400 ;
        RECT 122.800 151.700 165.200 152.300 ;
        RECT 122.800 151.600 123.600 151.700 ;
        RECT 150.000 151.600 150.800 151.700 ;
        RECT 164.400 151.600 165.200 151.700 ;
        RECT 12.400 150.300 13.200 150.400 ;
        RECT 26.800 150.300 27.600 150.400 ;
        RECT 12.400 149.700 27.600 150.300 ;
        RECT 12.400 149.600 13.200 149.700 ;
        RECT 26.800 149.600 27.600 149.700 ;
        RECT 33.200 150.300 34.000 150.400 ;
        RECT 52.400 150.300 53.200 150.400 ;
        RECT 33.200 149.700 53.200 150.300 ;
        RECT 33.200 149.600 34.000 149.700 ;
        RECT 52.400 149.600 53.200 149.700 ;
        RECT 73.200 150.300 74.000 150.400 ;
        RECT 82.800 150.300 83.600 150.400 ;
        RECT 94.000 150.300 94.800 150.400 ;
        RECT 73.200 149.700 94.800 150.300 ;
        RECT 73.200 149.600 74.000 149.700 ;
        RECT 82.800 149.600 83.600 149.700 ;
        RECT 94.000 149.600 94.800 149.700 ;
        RECT 118.000 150.300 118.800 150.400 ;
        RECT 126.000 150.300 126.800 150.400 ;
        RECT 137.200 150.300 138.000 150.400 ;
        RECT 118.000 149.700 138.000 150.300 ;
        RECT 118.000 149.600 118.800 149.700 ;
        RECT 126.000 149.600 126.800 149.700 ;
        RECT 137.200 149.600 138.000 149.700 ;
        RECT 138.800 150.300 139.600 150.400 ;
        RECT 142.000 150.300 142.800 150.400 ;
        RECT 145.200 150.300 146.000 150.400 ;
        RECT 138.800 149.700 146.000 150.300 ;
        RECT 138.800 149.600 139.600 149.700 ;
        RECT 142.000 149.600 142.800 149.700 ;
        RECT 145.200 149.600 146.000 149.700 ;
        RECT 154.800 150.300 155.600 150.400 ;
        RECT 166.000 150.300 166.800 150.400 ;
        RECT 154.800 149.700 166.800 150.300 ;
        RECT 154.800 149.600 155.600 149.700 ;
        RECT 166.000 149.600 166.800 149.700 ;
        RECT 172.400 150.300 173.200 150.400 ;
        RECT 180.400 150.300 181.200 150.400 ;
        RECT 172.400 149.700 181.200 150.300 ;
        RECT 172.400 149.600 173.200 149.700 ;
        RECT 180.400 149.600 181.200 149.700 ;
        RECT 68.400 148.300 69.200 148.400 ;
        RECT 71.600 148.300 72.400 148.400 ;
        RECT 68.400 147.700 72.400 148.300 ;
        RECT 68.400 147.600 69.200 147.700 ;
        RECT 71.600 147.600 72.400 147.700 ;
        RECT 81.200 148.300 82.000 148.400 ;
        RECT 86.000 148.300 86.800 148.400 ;
        RECT 81.200 147.700 86.800 148.300 ;
        RECT 81.200 147.600 82.000 147.700 ;
        RECT 86.000 147.600 86.800 147.700 ;
        RECT 106.800 148.300 107.600 148.400 ;
        RECT 116.400 148.300 117.200 148.400 ;
        RECT 129.200 148.300 130.000 148.400 ;
        RECT 140.400 148.300 141.200 148.400 ;
        RECT 106.800 147.700 141.200 148.300 ;
        RECT 106.800 147.600 107.600 147.700 ;
        RECT 116.400 147.600 117.200 147.700 ;
        RECT 129.200 147.600 130.000 147.700 ;
        RECT 140.400 147.600 141.200 147.700 ;
        RECT 143.600 148.300 144.400 148.400 ;
        RECT 154.800 148.300 155.600 148.400 ;
        RECT 143.600 147.700 155.600 148.300 ;
        RECT 143.600 147.600 144.400 147.700 ;
        RECT 154.800 147.600 155.600 147.700 ;
        RECT 31.600 146.300 32.400 146.400 ;
        RECT 44.400 146.300 45.200 146.400 ;
        RECT 49.200 146.300 50.000 146.400 ;
        RECT 31.600 145.700 50.000 146.300 ;
        RECT 31.600 145.600 32.400 145.700 ;
        RECT 44.400 145.600 45.200 145.700 ;
        RECT 49.200 145.600 50.000 145.700 ;
        RECT 132.400 146.300 133.200 146.400 ;
        RECT 143.600 146.300 144.400 146.400 ;
        RECT 156.400 146.300 157.200 146.400 ;
        RECT 132.400 145.700 157.200 146.300 ;
        RECT 132.400 145.600 133.200 145.700 ;
        RECT 143.600 145.600 144.400 145.700 ;
        RECT 156.400 145.600 157.200 145.700 ;
        RECT 9.200 144.300 10.000 144.400 ;
        RECT 20.400 144.300 21.200 144.400 ;
        RECT 30.000 144.300 30.800 144.400 ;
        RECT 46.000 144.300 46.800 144.400 ;
        RECT 9.200 143.700 46.800 144.300 ;
        RECT 9.200 143.600 10.000 143.700 ;
        RECT 20.400 143.600 21.200 143.700 ;
        RECT 30.000 143.600 30.800 143.700 ;
        RECT 46.000 143.600 46.800 143.700 ;
        RECT 54.000 144.300 54.800 144.400 ;
        RECT 65.200 144.300 66.000 144.400 ;
        RECT 54.000 143.700 66.000 144.300 ;
        RECT 54.000 143.600 54.800 143.700 ;
        RECT 65.200 143.600 66.000 143.700 ;
        RECT 137.200 144.300 138.000 144.400 ;
        RECT 143.600 144.300 144.400 144.400 ;
        RECT 137.200 143.700 144.400 144.300 ;
        RECT 137.200 143.600 138.000 143.700 ;
        RECT 143.600 143.600 144.400 143.700 ;
        RECT 174.000 142.300 174.800 142.400 ;
        RECT 193.200 142.300 194.000 142.400 ;
        RECT 174.000 141.700 194.000 142.300 ;
        RECT 174.000 141.600 174.800 141.700 ;
        RECT 193.200 141.600 194.000 141.700 ;
        RECT 62.000 138.300 62.800 138.400 ;
        RECT 84.400 138.300 85.200 138.400 ;
        RECT 62.000 137.700 85.200 138.300 ;
        RECT 62.000 137.600 62.800 137.700 ;
        RECT 84.400 137.600 85.200 137.700 ;
        RECT 142.000 138.300 142.800 138.400 ;
        RECT 146.800 138.300 147.600 138.400 ;
        RECT 142.000 137.700 147.600 138.300 ;
        RECT 142.000 137.600 142.800 137.700 ;
        RECT 146.800 137.600 147.600 137.700 ;
        RECT 15.600 136.300 16.400 136.400 ;
        RECT 20.400 136.300 21.200 136.400 ;
        RECT 15.600 135.700 21.200 136.300 ;
        RECT 15.600 135.600 16.400 135.700 ;
        RECT 20.400 135.600 21.200 135.700 ;
        RECT 25.200 136.300 26.000 136.400 ;
        RECT 34.800 136.300 35.600 136.400 ;
        RECT 25.200 135.700 35.600 136.300 ;
        RECT 25.200 135.600 26.000 135.700 ;
        RECT 34.800 135.600 35.600 135.700 ;
        RECT 47.600 136.300 48.400 136.400 ;
        RECT 50.800 136.300 51.600 136.400 ;
        RECT 63.600 136.300 64.400 136.400 ;
        RECT 47.600 135.700 64.400 136.300 ;
        RECT 47.600 135.600 48.400 135.700 ;
        RECT 50.800 135.600 51.600 135.700 ;
        RECT 63.600 135.600 64.400 135.700 ;
        RECT 119.600 136.300 120.400 136.400 ;
        RECT 122.800 136.300 123.600 136.400 ;
        RECT 119.600 135.700 123.600 136.300 ;
        RECT 119.600 135.600 120.400 135.700 ;
        RECT 122.800 135.600 123.600 135.700 ;
        RECT 145.200 136.300 146.000 136.400 ;
        RECT 150.000 136.300 150.800 136.400 ;
        RECT 145.200 135.700 150.800 136.300 ;
        RECT 145.200 135.600 146.000 135.700 ;
        RECT 150.000 135.600 150.800 135.700 ;
        RECT 156.400 136.300 157.200 136.400 ;
        RECT 161.200 136.300 162.000 136.400 ;
        RECT 156.400 135.700 162.000 136.300 ;
        RECT 156.400 135.600 157.200 135.700 ;
        RECT 161.200 135.600 162.000 135.700 ;
        RECT 23.600 134.300 24.400 134.400 ;
        RECT 26.800 134.300 27.600 134.400 ;
        RECT 23.600 133.700 27.600 134.300 ;
        RECT 23.600 133.600 24.400 133.700 ;
        RECT 26.800 133.600 27.600 133.700 ;
        RECT 28.400 134.300 29.200 134.400 ;
        RECT 44.400 134.300 45.200 134.400 ;
        RECT 28.400 133.700 45.200 134.300 ;
        RECT 28.400 133.600 29.200 133.700 ;
        RECT 44.400 133.600 45.200 133.700 ;
        RECT 100.400 134.300 101.200 134.400 ;
        RECT 110.000 134.300 110.800 134.400 ;
        RECT 100.400 133.700 110.800 134.300 ;
        RECT 100.400 133.600 101.200 133.700 ;
        RECT 110.000 133.600 110.800 133.700 ;
        RECT 137.200 134.300 138.000 134.400 ;
        RECT 153.200 134.300 154.000 134.400 ;
        RECT 159.600 134.300 160.400 134.400 ;
        RECT 137.200 133.700 160.400 134.300 ;
        RECT 137.200 133.600 138.000 133.700 ;
        RECT 153.200 133.600 154.000 133.700 ;
        RECT 159.600 133.600 160.400 133.700 ;
        RECT 166.000 134.300 166.800 134.400 ;
        RECT 172.400 134.300 173.200 134.400 ;
        RECT 166.000 133.700 173.200 134.300 ;
        RECT 166.000 133.600 166.800 133.700 ;
        RECT 172.400 133.600 173.200 133.700 ;
        RECT 1.200 132.300 2.000 132.400 ;
        RECT 4.400 132.300 5.200 132.400 ;
        RECT 10.800 132.300 11.600 132.400 ;
        RECT 15.600 132.300 16.400 132.400 ;
        RECT 58.800 132.300 59.600 132.400 ;
        RECT 1.200 131.700 59.600 132.300 ;
        RECT 1.200 131.600 2.000 131.700 ;
        RECT 4.400 131.600 5.200 131.700 ;
        RECT 10.800 131.600 11.600 131.700 ;
        RECT 15.600 131.600 16.400 131.700 ;
        RECT 58.800 131.600 59.600 131.700 ;
        RECT 63.600 132.300 64.400 132.400 ;
        RECT 73.200 132.300 74.000 132.400 ;
        RECT 63.600 131.700 74.000 132.300 ;
        RECT 63.600 131.600 64.400 131.700 ;
        RECT 73.200 131.600 74.000 131.700 ;
        RECT 79.600 132.300 80.400 132.400 ;
        RECT 95.600 132.300 96.400 132.400 ;
        RECT 79.600 131.700 96.400 132.300 ;
        RECT 79.600 131.600 80.400 131.700 ;
        RECT 95.600 131.600 96.400 131.700 ;
        RECT 114.800 132.300 115.600 132.400 ;
        RECT 122.800 132.300 123.600 132.400 ;
        RECT 114.800 131.700 123.600 132.300 ;
        RECT 114.800 131.600 115.600 131.700 ;
        RECT 122.800 131.600 123.600 131.700 ;
        RECT 130.800 132.300 131.600 132.400 ;
        RECT 135.600 132.300 136.400 132.400 ;
        RECT 151.600 132.300 152.400 132.400 ;
        RECT 156.400 132.300 157.200 132.400 ;
        RECT 130.800 131.700 157.200 132.300 ;
        RECT 130.800 131.600 131.600 131.700 ;
        RECT 135.600 131.600 136.400 131.700 ;
        RECT 151.600 131.600 152.400 131.700 ;
        RECT 156.400 131.600 157.200 131.700 ;
        RECT 12.400 130.300 13.200 130.400 ;
        RECT 18.800 130.300 19.600 130.400 ;
        RECT 36.400 130.300 37.200 130.400 ;
        RECT 12.400 129.700 37.200 130.300 ;
        RECT 12.400 129.600 13.200 129.700 ;
        RECT 18.800 129.600 19.600 129.700 ;
        RECT 36.400 129.600 37.200 129.700 ;
        RECT 68.400 130.300 69.200 130.400 ;
        RECT 84.400 130.300 85.200 130.400 ;
        RECT 68.400 129.700 85.200 130.300 ;
        RECT 68.400 129.600 69.200 129.700 ;
        RECT 84.400 129.600 85.200 129.700 ;
        RECT 103.600 130.300 104.400 130.400 ;
        RECT 127.600 130.300 128.400 130.400 ;
        RECT 132.400 130.300 133.200 130.400 ;
        RECT 103.600 129.700 133.200 130.300 ;
        RECT 103.600 129.600 104.400 129.700 ;
        RECT 127.600 129.600 128.400 129.700 ;
        RECT 132.400 129.600 133.200 129.700 ;
        RECT 159.600 130.300 160.400 130.400 ;
        RECT 167.600 130.300 168.400 130.400 ;
        RECT 159.600 129.700 168.400 130.300 ;
        RECT 159.600 129.600 160.400 129.700 ;
        RECT 167.600 129.600 168.400 129.700 ;
        RECT 36.400 128.300 37.200 128.400 ;
        RECT 57.200 128.300 58.000 128.400 ;
        RECT 36.400 127.700 58.000 128.300 ;
        RECT 36.400 127.600 37.200 127.700 ;
        RECT 57.200 127.600 58.000 127.700 ;
        RECT 60.400 128.300 61.200 128.400 ;
        RECT 63.600 128.300 64.400 128.400 ;
        RECT 71.600 128.300 72.400 128.400 ;
        RECT 78.000 128.300 78.800 128.400 ;
        RECT 87.600 128.300 88.400 128.400 ;
        RECT 60.400 127.700 88.400 128.300 ;
        RECT 60.400 127.600 61.200 127.700 ;
        RECT 63.600 127.600 64.400 127.700 ;
        RECT 71.600 127.600 72.400 127.700 ;
        RECT 78.000 127.600 78.800 127.700 ;
        RECT 87.600 127.600 88.400 127.700 ;
        RECT 126.000 128.300 126.800 128.400 ;
        RECT 130.800 128.300 131.600 128.400 ;
        RECT 126.000 127.700 131.600 128.300 ;
        RECT 126.000 127.600 126.800 127.700 ;
        RECT 130.800 127.600 131.600 127.700 ;
        RECT 138.800 128.300 139.600 128.400 ;
        RECT 177.200 128.300 178.000 128.400 ;
        RECT 138.800 127.700 178.000 128.300 ;
        RECT 138.800 127.600 139.600 127.700 ;
        RECT 177.200 127.600 178.000 127.700 ;
        RECT 46.000 126.300 46.800 126.400 ;
        RECT 65.200 126.300 66.000 126.400 ;
        RECT 46.000 125.700 66.000 126.300 ;
        RECT 46.000 125.600 46.800 125.700 ;
        RECT 65.200 125.600 66.000 125.700 ;
        RECT 38.000 124.300 38.800 124.400 ;
        RECT 46.000 124.300 46.800 124.400 ;
        RECT 79.600 124.300 80.400 124.400 ;
        RECT 38.000 123.700 80.400 124.300 ;
        RECT 38.000 123.600 38.800 123.700 ;
        RECT 46.000 123.600 46.800 123.700 ;
        RECT 79.600 123.600 80.400 123.700 ;
        RECT 97.200 124.300 98.000 124.400 ;
        RECT 98.800 124.300 99.600 124.400 ;
        RECT 97.200 123.700 99.600 124.300 ;
        RECT 97.200 123.600 98.000 123.700 ;
        RECT 98.800 123.600 99.600 123.700 ;
        RECT 41.200 118.300 42.000 118.400 ;
        RECT 119.600 118.300 120.400 118.400 ;
        RECT 41.200 117.700 120.400 118.300 ;
        RECT 41.200 117.600 42.000 117.700 ;
        RECT 119.600 117.600 120.400 117.700 ;
        RECT 122.800 118.300 123.600 118.400 ;
        RECT 146.800 118.300 147.600 118.400 ;
        RECT 122.800 117.700 147.600 118.300 ;
        RECT 122.800 117.600 123.600 117.700 ;
        RECT 146.800 117.600 147.600 117.700 ;
        RECT 38.000 114.300 38.800 114.400 ;
        RECT 47.600 114.300 48.400 114.400 ;
        RECT 58.800 114.300 59.600 114.400 ;
        RECT 116.400 114.300 117.200 114.400 ;
        RECT 38.000 113.700 117.200 114.300 ;
        RECT 38.000 113.600 38.800 113.700 ;
        RECT 47.600 113.600 48.400 113.700 ;
        RECT 58.800 113.600 59.600 113.700 ;
        RECT 116.400 113.600 117.200 113.700 ;
        RECT 119.600 114.300 120.400 114.400 ;
        RECT 129.200 114.300 130.000 114.400 ;
        RECT 119.600 113.700 130.000 114.300 ;
        RECT 119.600 113.600 120.400 113.700 ;
        RECT 129.200 113.600 130.000 113.700 ;
        RECT 18.800 112.300 19.600 112.400 ;
        RECT 25.200 112.300 26.000 112.400 ;
        RECT 18.800 111.700 26.000 112.300 ;
        RECT 18.800 111.600 19.600 111.700 ;
        RECT 25.200 111.600 26.000 111.700 ;
        RECT 47.600 112.300 48.400 112.400 ;
        RECT 50.800 112.300 51.600 112.400 ;
        RECT 63.600 112.300 64.400 112.400 ;
        RECT 47.600 111.700 64.400 112.300 ;
        RECT 47.600 111.600 48.400 111.700 ;
        RECT 50.800 111.600 51.600 111.700 ;
        RECT 63.600 111.600 64.400 111.700 ;
        RECT 70.000 112.300 70.800 112.400 ;
        RECT 73.200 112.300 74.000 112.400 ;
        RECT 70.000 111.700 74.000 112.300 ;
        RECT 70.000 111.600 70.800 111.700 ;
        RECT 73.200 111.600 74.000 111.700 ;
        RECT 92.400 112.300 93.200 112.400 ;
        RECT 111.600 112.300 112.400 112.400 ;
        RECT 92.400 111.700 112.400 112.300 ;
        RECT 92.400 111.600 93.200 111.700 ;
        RECT 111.600 111.600 112.400 111.700 ;
        RECT 126.000 112.300 126.800 112.400 ;
        RECT 129.200 112.300 130.000 112.400 ;
        RECT 126.000 111.700 130.000 112.300 ;
        RECT 126.000 111.600 126.800 111.700 ;
        RECT 129.200 111.600 130.000 111.700 ;
        RECT 154.800 112.300 155.600 112.400 ;
        RECT 167.600 112.300 168.400 112.400 ;
        RECT 170.800 112.300 171.600 112.400 ;
        RECT 154.800 111.700 171.600 112.300 ;
        RECT 154.800 111.600 155.600 111.700 ;
        RECT 167.600 111.600 168.400 111.700 ;
        RECT 170.800 111.600 171.600 111.700 ;
        RECT 4.400 110.300 5.200 110.400 ;
        RECT 6.000 110.300 6.800 110.400 ;
        RECT 28.400 110.300 29.200 110.400 ;
        RECT 4.400 109.700 29.200 110.300 ;
        RECT 4.400 109.600 5.200 109.700 ;
        RECT 6.000 109.600 6.800 109.700 ;
        RECT 28.400 109.600 29.200 109.700 ;
        RECT 60.400 110.300 61.200 110.400 ;
        RECT 65.200 110.300 66.000 110.400 ;
        RECT 60.400 109.700 66.000 110.300 ;
        RECT 60.400 109.600 61.200 109.700 ;
        RECT 65.200 109.600 66.000 109.700 ;
        RECT 73.200 110.300 74.000 110.400 ;
        RECT 82.800 110.300 83.600 110.400 ;
        RECT 87.600 110.300 88.400 110.400 ;
        RECT 94.000 110.300 94.800 110.400 ;
        RECT 73.200 109.700 94.800 110.300 ;
        RECT 73.200 109.600 74.000 109.700 ;
        RECT 82.800 109.600 83.600 109.700 ;
        RECT 87.600 109.600 88.400 109.700 ;
        RECT 94.000 109.600 94.800 109.700 ;
        RECT 110.000 110.300 110.800 110.400 ;
        RECT 126.000 110.300 126.800 110.400 ;
        RECT 110.000 109.700 126.800 110.300 ;
        RECT 110.000 109.600 110.800 109.700 ;
        RECT 126.000 109.600 126.800 109.700 ;
        RECT 156.400 110.300 157.200 110.400 ;
        RECT 164.400 110.300 165.200 110.400 ;
        RECT 156.400 109.700 165.200 110.300 ;
        RECT 156.400 109.600 157.200 109.700 ;
        RECT 164.400 109.600 165.200 109.700 ;
        RECT 22.000 108.300 22.800 108.400 ;
        RECT 30.000 108.300 30.800 108.400 ;
        RECT 44.400 108.300 45.200 108.400 ;
        RECT 49.200 108.300 50.000 108.400 ;
        RECT 22.000 107.700 50.000 108.300 ;
        RECT 22.000 107.600 22.800 107.700 ;
        RECT 30.000 107.600 30.800 107.700 ;
        RECT 44.400 107.600 45.200 107.700 ;
        RECT 49.200 107.600 50.000 107.700 ;
        RECT 89.200 108.300 90.000 108.400 ;
        RECT 95.600 108.300 96.400 108.400 ;
        RECT 89.200 107.700 96.400 108.300 ;
        RECT 89.200 107.600 90.000 107.700 ;
        RECT 95.600 107.600 96.400 107.700 ;
        RECT 111.600 108.300 112.400 108.400 ;
        RECT 146.800 108.300 147.600 108.400 ;
        RECT 162.800 108.300 163.600 108.400 ;
        RECT 111.600 107.700 163.600 108.300 ;
        RECT 111.600 107.600 112.400 107.700 ;
        RECT 146.800 107.600 147.600 107.700 ;
        RECT 162.800 107.600 163.600 107.700 ;
        RECT 164.400 108.300 165.200 108.400 ;
        RECT 174.000 108.300 174.800 108.400 ;
        RECT 188.400 108.300 189.200 108.400 ;
        RECT 164.400 107.700 189.200 108.300 ;
        RECT 164.400 107.600 165.200 107.700 ;
        RECT 174.000 107.600 174.800 107.700 ;
        RECT 188.400 107.600 189.200 107.700 ;
        RECT 34.800 106.300 35.600 106.400 ;
        RECT 39.600 106.300 40.400 106.400 ;
        RECT 34.800 105.700 40.400 106.300 ;
        RECT 34.800 105.600 35.600 105.700 ;
        RECT 39.600 105.600 40.400 105.700 ;
        RECT 86.000 106.300 86.800 106.400 ;
        RECT 90.800 106.300 91.600 106.400 ;
        RECT 86.000 105.700 91.600 106.300 ;
        RECT 86.000 105.600 86.800 105.700 ;
        RECT 90.800 105.600 91.600 105.700 ;
        RECT 126.000 106.300 126.800 106.400 ;
        RECT 143.600 106.300 144.400 106.400 ;
        RECT 126.000 105.700 144.400 106.300 ;
        RECT 126.000 105.600 126.800 105.700 ;
        RECT 143.600 105.600 144.400 105.700 ;
        RECT 188.400 106.300 189.200 106.400 ;
        RECT 193.200 106.300 194.000 106.400 ;
        RECT 188.400 105.700 194.000 106.300 ;
        RECT 188.400 105.600 189.200 105.700 ;
        RECT 193.200 105.600 194.000 105.700 ;
        RECT 74.800 104.300 75.600 104.400 ;
        RECT 79.600 104.300 80.400 104.400 ;
        RECT 84.400 104.300 85.200 104.400 ;
        RECT 74.800 103.700 85.200 104.300 ;
        RECT 74.800 103.600 75.600 103.700 ;
        RECT 79.600 103.600 80.400 103.700 ;
        RECT 84.400 103.600 85.200 103.700 ;
        RECT 122.800 104.300 123.600 104.400 ;
        RECT 126.000 104.300 126.800 104.400 ;
        RECT 122.800 103.700 126.800 104.300 ;
        RECT 122.800 103.600 123.600 103.700 ;
        RECT 126.000 103.600 126.800 103.700 ;
        RECT 145.200 104.300 146.000 104.400 ;
        RECT 172.400 104.300 173.200 104.400 ;
        RECT 145.200 103.700 173.200 104.300 ;
        RECT 145.200 103.600 146.000 103.700 ;
        RECT 172.400 103.600 173.200 103.700 ;
        RECT 63.600 102.300 64.400 102.400 ;
        RECT 121.200 102.300 122.000 102.400 ;
        RECT 63.600 101.700 122.000 102.300 ;
        RECT 63.600 101.600 64.400 101.700 ;
        RECT 121.200 101.600 122.000 101.700 ;
        RECT 142.000 102.300 142.800 102.400 ;
        RECT 180.400 102.300 181.200 102.400 ;
        RECT 142.000 101.700 181.200 102.300 ;
        RECT 142.000 101.600 142.800 101.700 ;
        RECT 180.400 101.600 181.200 101.700 ;
        RECT 143.600 100.300 144.400 100.400 ;
        RECT 170.800 100.300 171.600 100.400 ;
        RECT 183.600 100.300 184.400 100.400 ;
        RECT 191.600 100.300 192.400 100.400 ;
        RECT 143.600 99.700 192.400 100.300 ;
        RECT 143.600 99.600 144.400 99.700 ;
        RECT 170.800 99.600 171.600 99.700 ;
        RECT 183.600 99.600 184.400 99.700 ;
        RECT 191.600 99.600 192.400 99.700 ;
        RECT 41.200 98.300 42.000 98.400 ;
        RECT 46.000 98.300 46.800 98.400 ;
        RECT 41.200 97.700 46.800 98.300 ;
        RECT 41.200 97.600 42.000 97.700 ;
        RECT 46.000 97.600 46.800 97.700 ;
        RECT 68.400 98.300 69.200 98.400 ;
        RECT 84.400 98.300 85.200 98.400 ;
        RECT 89.200 98.300 90.000 98.400 ;
        RECT 68.400 97.700 90.000 98.300 ;
        RECT 68.400 97.600 69.200 97.700 ;
        RECT 84.400 97.600 85.200 97.700 ;
        RECT 89.200 97.600 90.000 97.700 ;
        RECT 137.200 98.300 138.000 98.400 ;
        RECT 159.600 98.300 160.400 98.400 ;
        RECT 169.200 98.300 170.000 98.400 ;
        RECT 188.400 98.300 189.200 98.400 ;
        RECT 137.200 97.700 189.200 98.300 ;
        RECT 137.200 97.600 138.000 97.700 ;
        RECT 159.600 97.600 160.400 97.700 ;
        RECT 169.200 97.600 170.000 97.700 ;
        RECT 188.400 97.600 189.200 97.700 ;
        RECT 12.400 96.300 13.200 96.400 ;
        RECT 25.200 96.300 26.000 96.400 ;
        RECT 12.400 95.700 26.000 96.300 ;
        RECT 12.400 95.600 13.200 95.700 ;
        RECT 25.200 95.600 26.000 95.700 ;
        RECT 63.600 96.300 64.400 96.400 ;
        RECT 70.000 96.300 70.800 96.400 ;
        RECT 63.600 95.700 70.800 96.300 ;
        RECT 63.600 95.600 64.400 95.700 ;
        RECT 70.000 95.600 70.800 95.700 ;
        RECT 82.800 96.300 83.600 96.400 ;
        RECT 87.600 96.300 88.400 96.400 ;
        RECT 82.800 95.700 88.400 96.300 ;
        RECT 82.800 95.600 83.600 95.700 ;
        RECT 87.600 95.600 88.400 95.700 ;
        RECT 114.800 96.300 115.600 96.400 ;
        RECT 145.200 96.300 146.000 96.400 ;
        RECT 114.800 95.700 146.000 96.300 ;
        RECT 114.800 95.600 115.600 95.700 ;
        RECT 145.200 95.600 146.000 95.700 ;
        RECT 148.400 96.300 149.200 96.400 ;
        RECT 153.200 96.300 154.000 96.400 ;
        RECT 148.400 95.700 154.000 96.300 ;
        RECT 148.400 95.600 149.200 95.700 ;
        RECT 153.200 95.600 154.000 95.700 ;
        RECT 18.800 94.300 19.600 94.400 ;
        RECT 31.600 94.300 32.400 94.400 ;
        RECT 18.800 93.700 32.400 94.300 ;
        RECT 18.800 93.600 19.600 93.700 ;
        RECT 31.600 93.600 32.400 93.700 ;
        RECT 58.800 94.300 59.600 94.400 ;
        RECT 70.000 94.300 70.800 94.400 ;
        RECT 58.800 93.700 70.800 94.300 ;
        RECT 58.800 93.600 59.600 93.700 ;
        RECT 70.000 93.600 70.800 93.700 ;
        RECT 114.800 94.300 115.600 94.400 ;
        RECT 121.200 94.300 122.000 94.400 ;
        RECT 114.800 93.700 122.000 94.300 ;
        RECT 114.800 93.600 115.600 93.700 ;
        RECT 121.200 93.600 122.000 93.700 ;
        RECT 129.200 94.300 130.000 94.400 ;
        RECT 134.000 94.300 134.800 94.400 ;
        RECT 143.600 94.300 144.400 94.400 ;
        RECT 129.200 93.700 144.400 94.300 ;
        RECT 129.200 93.600 130.000 93.700 ;
        RECT 134.000 93.600 134.800 93.700 ;
        RECT 143.600 93.600 144.400 93.700 ;
        RECT 145.200 94.300 146.000 94.400 ;
        RECT 151.600 94.300 152.400 94.400 ;
        RECT 158.000 94.300 158.800 94.400 ;
        RECT 166.000 94.300 166.800 94.400 ;
        RECT 145.200 93.700 166.800 94.300 ;
        RECT 145.200 93.600 146.000 93.700 ;
        RECT 151.600 93.600 152.400 93.700 ;
        RECT 158.000 93.600 158.800 93.700 ;
        RECT 166.000 93.600 166.800 93.700 ;
        RECT 9.200 92.300 10.000 92.400 ;
        RECT 36.400 92.300 37.200 92.400 ;
        RECT 41.200 92.300 42.000 92.400 ;
        RECT 9.200 91.700 42.000 92.300 ;
        RECT 9.200 91.600 10.000 91.700 ;
        RECT 36.400 91.600 37.200 91.700 ;
        RECT 41.200 91.600 42.000 91.700 ;
        RECT 44.400 92.300 45.200 92.400 ;
        RECT 60.400 92.300 61.200 92.400 ;
        RECT 44.400 91.700 61.200 92.300 ;
        RECT 44.400 91.600 45.200 91.700 ;
        RECT 60.400 91.600 61.200 91.700 ;
        RECT 76.400 92.300 77.200 92.400 ;
        RECT 79.600 92.300 80.400 92.400 ;
        RECT 76.400 91.700 80.400 92.300 ;
        RECT 76.400 91.600 77.200 91.700 ;
        RECT 79.600 91.600 80.400 91.700 ;
        RECT 87.600 92.300 88.400 92.400 ;
        RECT 98.800 92.300 99.600 92.400 ;
        RECT 87.600 91.700 99.600 92.300 ;
        RECT 87.600 91.600 88.400 91.700 ;
        RECT 98.800 91.600 99.600 91.700 ;
        RECT 119.600 92.300 120.400 92.400 ;
        RECT 126.000 92.300 126.800 92.400 ;
        RECT 119.600 91.700 126.800 92.300 ;
        RECT 119.600 91.600 120.400 91.700 ;
        RECT 126.000 91.600 126.800 91.700 ;
        RECT 130.800 92.300 131.600 92.400 ;
        RECT 137.200 92.300 138.000 92.400 ;
        RECT 130.800 91.700 138.000 92.300 ;
        RECT 130.800 91.600 131.600 91.700 ;
        RECT 137.200 91.600 138.000 91.700 ;
        RECT 150.000 92.300 150.800 92.400 ;
        RECT 156.400 92.300 157.200 92.400 ;
        RECT 164.400 92.300 165.200 92.400 ;
        RECT 150.000 91.700 165.200 92.300 ;
        RECT 150.000 91.600 150.800 91.700 ;
        RECT 156.400 91.600 157.200 91.700 ;
        RECT 164.400 91.600 165.200 91.700 ;
        RECT 54.000 90.300 54.800 90.400 ;
        RECT 73.200 90.300 74.000 90.400 ;
        RECT 78.000 90.300 78.800 90.400 ;
        RECT 89.200 90.300 90.000 90.400 ;
        RECT 108.400 90.300 109.200 90.400 ;
        RECT 54.000 89.700 109.200 90.300 ;
        RECT 54.000 89.600 54.800 89.700 ;
        RECT 73.200 89.600 74.000 89.700 ;
        RECT 78.000 89.600 78.800 89.700 ;
        RECT 89.200 89.600 90.000 89.700 ;
        RECT 108.400 89.600 109.200 89.700 ;
        RECT 30.000 84.300 30.800 84.400 ;
        RECT 36.400 84.300 37.200 84.400 ;
        RECT 30.000 83.700 37.200 84.300 ;
        RECT 30.000 83.600 30.800 83.700 ;
        RECT 36.400 83.600 37.200 83.700 ;
        RECT 26.800 82.300 27.600 82.400 ;
        RECT 30.000 82.300 30.800 82.400 ;
        RECT 26.800 81.700 30.800 82.300 ;
        RECT 26.800 81.600 27.600 81.700 ;
        RECT 30.000 81.600 30.800 81.700 ;
        RECT 86.000 82.300 86.800 82.400 ;
        RECT 95.600 82.300 96.400 82.400 ;
        RECT 108.400 82.300 109.200 82.400 ;
        RECT 86.000 81.700 109.200 82.300 ;
        RECT 86.000 81.600 86.800 81.700 ;
        RECT 95.600 81.600 96.400 81.700 ;
        RECT 108.400 81.600 109.200 81.700 ;
        RECT 122.800 80.300 123.600 80.400 ;
        RECT 127.600 80.300 128.400 80.400 ;
        RECT 132.400 80.300 133.200 80.400 ;
        RECT 122.800 79.700 133.200 80.300 ;
        RECT 122.800 79.600 123.600 79.700 ;
        RECT 127.600 79.600 128.400 79.700 ;
        RECT 132.400 79.600 133.200 79.700 ;
        RECT 68.400 78.300 69.200 78.400 ;
        RECT 73.200 78.300 74.000 78.400 ;
        RECT 68.400 77.700 74.000 78.300 ;
        RECT 68.400 77.600 69.200 77.700 ;
        RECT 73.200 77.600 74.000 77.700 ;
        RECT 153.200 74.300 154.000 74.400 ;
        RECT 178.800 74.300 179.600 74.400 ;
        RECT 153.200 73.700 179.600 74.300 ;
        RECT 153.200 73.600 154.000 73.700 ;
        RECT 178.800 73.600 179.600 73.700 ;
        RECT 10.800 72.300 11.600 72.400 ;
        RECT 14.000 72.300 14.800 72.400 ;
        RECT 10.800 71.700 14.800 72.300 ;
        RECT 10.800 71.600 11.600 71.700 ;
        RECT 14.000 71.600 14.800 71.700 ;
        RECT 17.200 72.300 18.000 72.400 ;
        RECT 20.400 72.300 21.200 72.400 ;
        RECT 17.200 71.700 21.200 72.300 ;
        RECT 17.200 71.600 18.000 71.700 ;
        RECT 20.400 71.600 21.200 71.700 ;
        RECT 39.600 72.300 40.400 72.400 ;
        RECT 47.600 72.300 48.400 72.400 ;
        RECT 39.600 71.700 48.400 72.300 ;
        RECT 39.600 71.600 40.400 71.700 ;
        RECT 47.600 71.600 48.400 71.700 ;
        RECT 134.000 72.300 134.800 72.400 ;
        RECT 146.800 72.300 147.600 72.400 ;
        RECT 134.000 71.700 147.600 72.300 ;
        RECT 134.000 71.600 134.800 71.700 ;
        RECT 146.800 71.600 147.600 71.700 ;
        RECT 4.400 70.300 5.200 70.400 ;
        RECT 9.200 70.300 10.000 70.400 ;
        RECT 23.600 70.300 24.400 70.400 ;
        RECT 31.600 70.300 32.400 70.400 ;
        RECT 60.400 70.300 61.200 70.400 ;
        RECT 4.400 69.700 61.200 70.300 ;
        RECT 4.400 69.600 5.200 69.700 ;
        RECT 9.200 69.600 10.000 69.700 ;
        RECT 23.600 69.600 24.400 69.700 ;
        RECT 31.600 69.600 32.400 69.700 ;
        RECT 60.400 69.600 61.200 69.700 ;
        RECT 98.800 70.300 99.600 70.400 ;
        RECT 105.200 70.300 106.000 70.400 ;
        RECT 127.600 70.300 128.400 70.400 ;
        RECT 98.800 69.700 128.400 70.300 ;
        RECT 98.800 69.600 99.600 69.700 ;
        RECT 105.200 69.600 106.000 69.700 ;
        RECT 127.600 69.600 128.400 69.700 ;
        RECT 138.800 70.300 139.600 70.400 ;
        RECT 142.000 70.300 142.800 70.400 ;
        RECT 138.800 69.700 142.800 70.300 ;
        RECT 138.800 69.600 139.600 69.700 ;
        RECT 142.000 69.600 142.800 69.700 ;
        RECT 145.200 70.300 146.000 70.400 ;
        RECT 166.000 70.300 166.800 70.400 ;
        RECT 145.200 69.700 166.800 70.300 ;
        RECT 145.200 69.600 146.000 69.700 ;
        RECT 166.000 69.600 166.800 69.700 ;
        RECT 30.000 68.300 30.800 68.400 ;
        RECT 38.000 68.300 38.800 68.400 ;
        RECT 30.000 67.700 38.800 68.300 ;
        RECT 30.000 67.600 30.800 67.700 ;
        RECT 38.000 67.600 38.800 67.700 ;
        RECT 102.000 68.300 102.800 68.400 ;
        RECT 111.600 68.300 112.400 68.400 ;
        RECT 102.000 67.700 112.400 68.300 ;
        RECT 102.000 67.600 102.800 67.700 ;
        RECT 111.600 67.600 112.400 67.700 ;
        RECT 22.000 66.300 22.800 66.400 ;
        RECT 26.800 66.300 27.600 66.400 ;
        RECT 30.000 66.300 30.800 66.400 ;
        RECT 33.200 66.300 34.000 66.400 ;
        RECT 22.000 65.700 34.000 66.300 ;
        RECT 22.000 65.600 22.800 65.700 ;
        RECT 26.800 65.600 27.600 65.700 ;
        RECT 30.000 65.600 30.800 65.700 ;
        RECT 33.200 65.600 34.000 65.700 ;
        RECT 38.000 66.300 38.800 66.400 ;
        RECT 41.200 66.300 42.000 66.400 ;
        RECT 38.000 65.700 42.000 66.300 ;
        RECT 38.000 65.600 38.800 65.700 ;
        RECT 41.200 65.600 42.000 65.700 ;
        RECT 95.600 66.300 96.400 66.400 ;
        RECT 100.400 66.300 101.200 66.400 ;
        RECT 95.600 65.700 101.200 66.300 ;
        RECT 95.600 65.600 96.400 65.700 ;
        RECT 100.400 65.600 101.200 65.700 ;
        RECT 126.000 66.300 126.800 66.400 ;
        RECT 151.600 66.300 152.400 66.400 ;
        RECT 126.000 65.700 152.400 66.300 ;
        RECT 126.000 65.600 126.800 65.700 ;
        RECT 151.600 65.600 152.400 65.700 ;
        RECT 97.200 64.300 98.000 64.400 ;
        RECT 105.200 64.300 106.000 64.400 ;
        RECT 129.200 64.300 130.000 64.400 ;
        RECT 130.800 64.300 131.600 64.400 ;
        RECT 97.200 63.700 131.600 64.300 ;
        RECT 97.200 63.600 98.000 63.700 ;
        RECT 105.200 63.600 106.000 63.700 ;
        RECT 129.200 63.600 130.000 63.700 ;
        RECT 130.800 63.600 131.600 63.700 ;
        RECT 150.000 64.300 150.800 64.400 ;
        RECT 154.800 64.300 155.600 64.400 ;
        RECT 150.000 63.700 155.600 64.300 ;
        RECT 150.000 63.600 150.800 63.700 ;
        RECT 154.800 63.600 155.600 63.700 ;
        RECT 159.600 62.300 160.400 62.400 ;
        RECT 167.600 62.300 168.400 62.400 ;
        RECT 175.600 62.300 176.400 62.400 ;
        RECT 159.600 61.700 176.400 62.300 ;
        RECT 159.600 61.600 160.400 61.700 ;
        RECT 167.600 61.600 168.400 61.700 ;
        RECT 175.600 61.600 176.400 61.700 ;
        RECT 153.200 60.300 154.000 60.400 ;
        RECT 169.200 60.300 170.000 60.400 ;
        RECT 153.200 59.700 170.000 60.300 ;
        RECT 153.200 59.600 154.000 59.700 ;
        RECT 169.200 59.600 170.000 59.700 ;
        RECT 6.000 58.300 6.800 58.400 ;
        RECT 14.000 58.300 14.800 58.400 ;
        RECT 26.800 58.300 27.600 58.400 ;
        RECT 6.000 57.700 27.600 58.300 ;
        RECT 6.000 57.600 6.800 57.700 ;
        RECT 14.000 57.600 14.800 57.700 ;
        RECT 26.800 57.600 27.600 57.700 ;
        RECT 127.600 58.300 128.400 58.400 ;
        RECT 145.200 58.300 146.000 58.400 ;
        RECT 127.600 57.700 146.000 58.300 ;
        RECT 127.600 57.600 128.400 57.700 ;
        RECT 145.200 57.600 146.000 57.700 ;
        RECT 146.800 58.300 147.600 58.400 ;
        RECT 174.000 58.300 174.800 58.400 ;
        RECT 146.800 57.700 174.800 58.300 ;
        RECT 146.800 57.600 147.600 57.700 ;
        RECT 174.000 57.600 174.800 57.700 ;
        RECT 89.200 56.300 90.000 56.400 ;
        RECT 110.000 56.300 110.800 56.400 ;
        RECT 89.200 55.700 110.800 56.300 ;
        RECT 89.200 55.600 90.000 55.700 ;
        RECT 110.000 55.600 110.800 55.700 ;
        RECT 138.800 56.300 139.600 56.400 ;
        RECT 142.000 56.300 142.800 56.400 ;
        RECT 138.800 55.700 142.800 56.300 ;
        RECT 138.800 55.600 139.600 55.700 ;
        RECT 142.000 55.600 142.800 55.700 ;
        RECT 143.600 56.300 144.400 56.400 ;
        RECT 158.000 56.300 158.800 56.400 ;
        RECT 143.600 55.700 158.800 56.300 ;
        RECT 143.600 55.600 144.400 55.700 ;
        RECT 158.000 55.600 158.800 55.700 ;
        RECT 172.400 56.300 173.200 56.400 ;
        RECT 180.400 56.300 181.200 56.400 ;
        RECT 172.400 55.700 181.200 56.300 ;
        RECT 172.400 55.600 173.200 55.700 ;
        RECT 180.400 55.600 181.200 55.700 ;
        RECT 22.000 54.300 22.800 54.400 ;
        RECT 31.600 54.300 32.400 54.400 ;
        RECT 47.600 54.300 48.400 54.400 ;
        RECT 52.400 54.300 53.200 54.400 ;
        RECT 22.000 53.700 53.200 54.300 ;
        RECT 22.000 53.600 22.800 53.700 ;
        RECT 31.600 53.600 32.400 53.700 ;
        RECT 47.600 53.600 48.400 53.700 ;
        RECT 52.400 53.600 53.200 53.700 ;
        RECT 116.400 54.300 117.200 54.400 ;
        RECT 158.000 54.300 158.800 54.400 ;
        RECT 166.000 54.300 166.800 54.400 ;
        RECT 116.400 53.700 166.800 54.300 ;
        RECT 116.400 53.600 117.200 53.700 ;
        RECT 158.000 53.600 158.800 53.700 ;
        RECT 166.000 53.600 166.800 53.700 ;
        RECT 180.400 54.300 181.200 54.400 ;
        RECT 183.600 54.300 184.400 54.400 ;
        RECT 180.400 53.700 184.400 54.300 ;
        RECT 180.400 53.600 181.200 53.700 ;
        RECT 183.600 53.600 184.400 53.700 ;
        RECT 57.200 52.300 58.000 52.400 ;
        RECT 73.200 52.300 74.000 52.400 ;
        RECT 57.200 51.700 74.000 52.300 ;
        RECT 57.200 51.600 58.000 51.700 ;
        RECT 73.200 51.600 74.000 51.700 ;
        RECT 81.200 52.300 82.000 52.400 ;
        RECT 86.000 52.300 86.800 52.400 ;
        RECT 81.200 51.700 86.800 52.300 ;
        RECT 81.200 51.600 82.000 51.700 ;
        RECT 86.000 51.600 86.800 51.700 ;
        RECT 116.400 52.300 117.200 52.400 ;
        RECT 122.800 52.300 123.600 52.400 ;
        RECT 116.400 51.700 123.600 52.300 ;
        RECT 116.400 51.600 117.200 51.700 ;
        RECT 122.800 51.600 123.600 51.700 ;
        RECT 153.200 52.300 154.000 52.400 ;
        RECT 178.800 52.300 179.600 52.400 ;
        RECT 190.000 52.300 190.800 52.400 ;
        RECT 153.200 51.700 190.800 52.300 ;
        RECT 153.200 51.600 154.000 51.700 ;
        RECT 178.800 51.600 179.600 51.700 ;
        RECT 190.000 51.600 190.800 51.700 ;
        RECT 94.000 50.300 94.800 50.400 ;
        RECT 132.400 50.300 133.200 50.400 ;
        RECT 142.000 50.300 142.800 50.400 ;
        RECT 94.000 49.700 142.800 50.300 ;
        RECT 94.000 49.600 94.800 49.700 ;
        RECT 132.400 49.600 133.200 49.700 ;
        RECT 142.000 49.600 142.800 49.700 ;
        RECT 148.400 50.300 149.200 50.400 ;
        RECT 154.800 50.300 155.600 50.400 ;
        RECT 148.400 49.700 155.600 50.300 ;
        RECT 148.400 49.600 149.200 49.700 ;
        RECT 154.800 49.600 155.600 49.700 ;
        RECT 84.400 48.300 85.200 48.400 ;
        RECT 105.200 48.300 106.000 48.400 ;
        RECT 158.000 48.300 158.800 48.400 ;
        RECT 164.400 48.300 165.200 48.400 ;
        RECT 84.400 47.700 165.200 48.300 ;
        RECT 84.400 47.600 85.200 47.700 ;
        RECT 105.200 47.600 106.000 47.700 ;
        RECT 158.000 47.600 158.800 47.700 ;
        RECT 164.400 47.600 165.200 47.700 ;
        RECT 118.000 46.300 118.800 46.400 ;
        RECT 122.800 46.300 123.600 46.400 ;
        RECT 118.000 45.700 123.600 46.300 ;
        RECT 118.000 45.600 118.800 45.700 ;
        RECT 122.800 45.600 123.600 45.700 ;
        RECT 68.400 44.300 69.200 44.400 ;
        RECT 81.200 44.300 82.000 44.400 ;
        RECT 68.400 43.700 82.000 44.300 ;
        RECT 68.400 43.600 69.200 43.700 ;
        RECT 81.200 43.600 82.000 43.700 ;
        RECT 183.600 38.300 184.400 38.400 ;
        RECT 190.000 38.300 190.800 38.400 ;
        RECT 183.600 37.700 190.800 38.300 ;
        RECT 183.600 37.600 184.400 37.700 ;
        RECT 190.000 37.600 190.800 37.700 ;
        RECT 20.400 36.300 21.200 36.400 ;
        RECT 31.600 36.300 32.400 36.400 ;
        RECT 42.800 36.300 43.600 36.400 ;
        RECT 70.000 36.300 70.800 36.400 ;
        RECT 20.400 35.700 70.800 36.300 ;
        RECT 20.400 35.600 21.200 35.700 ;
        RECT 31.600 35.600 32.400 35.700 ;
        RECT 42.800 35.600 43.600 35.700 ;
        RECT 70.000 35.600 70.800 35.700 ;
        RECT 68.400 34.300 69.200 34.400 ;
        RECT 71.600 34.300 72.400 34.400 ;
        RECT 68.400 33.700 72.400 34.300 ;
        RECT 68.400 33.600 69.200 33.700 ;
        RECT 71.600 33.600 72.400 33.700 ;
        RECT 44.400 32.300 45.200 32.400 ;
        RECT 58.800 32.300 59.600 32.400 ;
        RECT 65.200 32.300 66.000 32.400 ;
        RECT 71.600 32.300 72.400 32.400 ;
        RECT 44.400 31.700 72.400 32.300 ;
        RECT 44.400 31.600 45.200 31.700 ;
        RECT 58.800 31.600 59.600 31.700 ;
        RECT 65.200 31.600 66.000 31.700 ;
        RECT 71.600 31.600 72.400 31.700 ;
        RECT 73.200 32.300 74.000 32.400 ;
        RECT 98.800 32.300 99.600 32.400 ;
        RECT 73.200 31.700 99.600 32.300 ;
        RECT 73.200 31.600 74.000 31.700 ;
        RECT 98.800 31.600 99.600 31.700 ;
        RECT 102.000 32.300 102.800 32.400 ;
        RECT 103.600 32.300 104.400 32.400 ;
        RECT 102.000 31.700 104.400 32.300 ;
        RECT 102.000 31.600 102.800 31.700 ;
        RECT 103.600 31.600 104.400 31.700 ;
        RECT 14.000 30.300 14.800 30.400 ;
        RECT 25.200 30.300 26.000 30.400 ;
        RECT 14.000 29.700 26.000 30.300 ;
        RECT 14.000 29.600 14.800 29.700 ;
        RECT 25.200 29.600 26.000 29.700 ;
        RECT 46.000 30.300 46.800 30.400 ;
        RECT 52.400 30.300 53.200 30.400 ;
        RECT 46.000 29.700 53.200 30.300 ;
        RECT 46.000 29.600 46.800 29.700 ;
        RECT 52.400 29.600 53.200 29.700 ;
        RECT 79.600 30.300 80.400 30.400 ;
        RECT 82.800 30.300 83.600 30.400 ;
        RECT 89.200 30.300 90.000 30.400 ;
        RECT 79.600 29.700 90.000 30.300 ;
        RECT 79.600 29.600 80.400 29.700 ;
        RECT 82.800 29.600 83.600 29.700 ;
        RECT 89.200 29.600 90.000 29.700 ;
        RECT 102.000 30.300 102.800 30.400 ;
        RECT 108.400 30.300 109.200 30.400 ;
        RECT 102.000 29.700 109.200 30.300 ;
        RECT 102.000 29.600 102.800 29.700 ;
        RECT 108.400 29.600 109.200 29.700 ;
        RECT 113.200 30.300 114.000 30.400 ;
        RECT 119.600 30.300 120.400 30.400 ;
        RECT 113.200 29.700 120.400 30.300 ;
        RECT 113.200 29.600 114.000 29.700 ;
        RECT 119.600 29.600 120.400 29.700 ;
        RECT 132.400 30.300 133.200 30.400 ;
        RECT 138.800 30.300 139.600 30.400 ;
        RECT 132.400 29.700 139.600 30.300 ;
        RECT 132.400 29.600 133.200 29.700 ;
        RECT 138.800 29.600 139.600 29.700 ;
        RECT 142.000 30.300 142.800 30.400 ;
        RECT 159.600 30.300 160.400 30.400 ;
        RECT 142.000 29.700 160.400 30.300 ;
        RECT 142.000 29.600 142.800 29.700 ;
        RECT 159.600 29.600 160.400 29.700 ;
        RECT 166.000 30.300 166.800 30.400 ;
        RECT 180.400 30.300 181.200 30.400 ;
        RECT 166.000 29.700 181.200 30.300 ;
        RECT 166.000 29.600 166.800 29.700 ;
        RECT 180.400 29.600 181.200 29.700 ;
        RECT 23.600 28.300 24.400 28.400 ;
        RECT 26.800 28.300 27.600 28.400 ;
        RECT 23.600 27.700 27.600 28.300 ;
        RECT 23.600 27.600 24.400 27.700 ;
        RECT 26.800 27.600 27.600 27.700 ;
        RECT 41.200 28.300 42.000 28.400 ;
        RECT 47.600 28.300 48.400 28.400 ;
        RECT 41.200 27.700 48.400 28.300 ;
        RECT 41.200 27.600 42.000 27.700 ;
        RECT 47.600 27.600 48.400 27.700 ;
        RECT 58.800 28.300 59.600 28.400 ;
        RECT 84.400 28.300 85.200 28.400 ;
        RECT 90.800 28.300 91.600 28.400 ;
        RECT 58.800 27.700 91.600 28.300 ;
        RECT 58.800 27.600 59.600 27.700 ;
        RECT 84.400 27.600 85.200 27.700 ;
        RECT 90.800 27.600 91.600 27.700 ;
        RECT 98.800 28.300 99.600 28.400 ;
        RECT 103.600 28.300 104.400 28.400 ;
        RECT 113.200 28.300 114.000 28.400 ;
        RECT 98.800 27.700 114.000 28.300 ;
        RECT 98.800 27.600 99.600 27.700 ;
        RECT 103.600 27.600 104.400 27.700 ;
        RECT 113.200 27.600 114.000 27.700 ;
        RECT 116.400 28.300 117.200 28.400 ;
        RECT 122.800 28.300 123.600 28.400 ;
        RECT 116.400 27.700 123.600 28.300 ;
        RECT 116.400 27.600 117.200 27.700 ;
        RECT 122.800 27.600 123.600 27.700 ;
        RECT 151.600 28.300 152.400 28.400 ;
        RECT 154.800 28.300 155.600 28.400 ;
        RECT 151.600 27.700 155.600 28.300 ;
        RECT 151.600 27.600 152.400 27.700 ;
        RECT 154.800 27.600 155.600 27.700 ;
        RECT 178.800 28.300 179.600 28.400 ;
        RECT 188.400 28.300 189.200 28.400 ;
        RECT 178.800 27.700 189.200 28.300 ;
        RECT 178.800 27.600 179.600 27.700 ;
        RECT 188.400 27.600 189.200 27.700 ;
        RECT 25.200 26.300 26.000 26.400 ;
        RECT 30.000 26.300 30.800 26.400 ;
        RECT 25.200 25.700 30.800 26.300 ;
        RECT 25.200 25.600 26.000 25.700 ;
        RECT 30.000 25.600 30.800 25.700 ;
        RECT 38.000 26.300 38.800 26.400 ;
        RECT 73.200 26.300 74.000 26.400 ;
        RECT 38.000 25.700 74.000 26.300 ;
        RECT 38.000 25.600 38.800 25.700 ;
        RECT 73.200 25.600 74.000 25.700 ;
        RECT 87.600 26.300 88.400 26.400 ;
        RECT 92.400 26.300 93.200 26.400 ;
        RECT 87.600 25.700 93.200 26.300 ;
        RECT 87.600 25.600 88.400 25.700 ;
        RECT 92.400 25.600 93.200 25.700 ;
        RECT 97.200 26.300 98.000 26.400 ;
        RECT 106.800 26.300 107.600 26.400 ;
        RECT 97.200 25.700 107.600 26.300 ;
        RECT 97.200 25.600 98.000 25.700 ;
        RECT 106.800 25.600 107.600 25.700 ;
        RECT 129.200 26.300 130.000 26.400 ;
        RECT 186.800 26.300 187.600 26.400 ;
        RECT 129.200 25.700 187.600 26.300 ;
        RECT 129.200 25.600 130.000 25.700 ;
        RECT 186.800 25.600 187.600 25.700 ;
        RECT 1.200 24.300 2.000 24.400 ;
        RECT 4.400 24.300 5.200 24.400 ;
        RECT 36.400 24.300 37.200 24.400 ;
        RECT 1.200 23.700 37.200 24.300 ;
        RECT 1.200 23.600 2.000 23.700 ;
        RECT 4.400 23.600 5.200 23.700 ;
        RECT 36.400 23.600 37.200 23.700 ;
        RECT 20.400 20.300 21.200 20.400 ;
        RECT 25.200 20.300 26.000 20.400 ;
        RECT 20.400 19.700 26.000 20.300 ;
        RECT 20.400 19.600 21.200 19.700 ;
        RECT 25.200 19.600 26.000 19.700 ;
        RECT 6.000 18.300 6.800 18.400 ;
        RECT 30.000 18.300 30.800 18.400 ;
        RECT 6.000 17.700 30.800 18.300 ;
        RECT 6.000 17.600 6.800 17.700 ;
        RECT 30.000 17.600 30.800 17.700 ;
        RECT 42.800 18.300 43.600 18.400 ;
        RECT 47.600 18.300 48.400 18.400 ;
        RECT 42.800 17.700 48.400 18.300 ;
        RECT 42.800 17.600 43.600 17.700 ;
        RECT 47.600 17.600 48.400 17.700 ;
        RECT 89.200 18.300 90.000 18.400 ;
        RECT 92.400 18.300 93.200 18.400 ;
        RECT 97.200 18.300 98.000 18.400 ;
        RECT 89.200 17.700 98.000 18.300 ;
        RECT 89.200 17.600 90.000 17.700 ;
        RECT 92.400 17.600 93.200 17.700 ;
        RECT 97.200 17.600 98.000 17.700 ;
        RECT 116.400 18.300 117.200 18.400 ;
        RECT 138.800 18.300 139.600 18.400 ;
        RECT 116.400 17.700 139.600 18.300 ;
        RECT 116.400 17.600 117.200 17.700 ;
        RECT 138.800 17.600 139.600 17.700 ;
        RECT 30.000 16.300 30.800 16.400 ;
        RECT 39.600 16.300 40.400 16.400 ;
        RECT 63.600 16.300 64.400 16.400 ;
        RECT 30.000 15.700 64.400 16.300 ;
        RECT 30.000 15.600 30.800 15.700 ;
        RECT 39.600 15.600 40.400 15.700 ;
        RECT 63.600 15.600 64.400 15.700 ;
        RECT 103.600 16.300 104.400 16.400 ;
        RECT 106.800 16.300 107.600 16.400 ;
        RECT 122.800 16.300 123.600 16.400 ;
        RECT 142.000 16.300 142.800 16.400 ;
        RECT 103.600 15.700 142.800 16.300 ;
        RECT 103.600 15.600 104.400 15.700 ;
        RECT 106.800 15.600 107.600 15.700 ;
        RECT 122.800 15.600 123.600 15.700 ;
        RECT 142.000 15.600 142.800 15.700 ;
        RECT 159.600 16.300 160.400 16.400 ;
        RECT 164.400 16.300 165.200 16.400 ;
        RECT 159.600 15.700 165.200 16.300 ;
        RECT 159.600 15.600 160.400 15.700 ;
        RECT 164.400 15.600 165.200 15.700 ;
        RECT 167.600 16.300 168.400 16.400 ;
        RECT 174.000 16.300 174.800 16.400 ;
        RECT 167.600 15.700 174.800 16.300 ;
        RECT 167.600 15.600 168.400 15.700 ;
        RECT 174.000 15.600 174.800 15.700 ;
        RECT 182.000 16.300 182.800 16.400 ;
        RECT 190.000 16.300 190.800 16.400 ;
        RECT 182.000 15.700 190.800 16.300 ;
        RECT 182.000 15.600 182.800 15.700 ;
        RECT 190.000 15.600 190.800 15.700 ;
        RECT 17.200 14.300 18.000 14.400 ;
        RECT 55.600 14.300 56.400 14.400 ;
        RECT 17.200 13.700 56.400 14.300 ;
        RECT 17.200 13.600 18.000 13.700 ;
        RECT 55.600 13.600 56.400 13.700 ;
        RECT 71.600 14.300 72.400 14.400 ;
        RECT 78.000 14.300 78.800 14.400 ;
        RECT 71.600 13.700 78.800 14.300 ;
        RECT 71.600 13.600 72.400 13.700 ;
        RECT 78.000 13.600 78.800 13.700 ;
        RECT 82.800 14.300 83.600 14.400 ;
        RECT 84.400 14.300 85.200 14.400 ;
        RECT 82.800 13.700 85.200 14.300 ;
        RECT 82.800 13.600 83.600 13.700 ;
        RECT 84.400 13.600 85.200 13.700 ;
        RECT 86.000 14.300 86.800 14.400 ;
        RECT 108.400 14.300 109.200 14.400 ;
        RECT 86.000 13.700 109.200 14.300 ;
        RECT 86.000 13.600 86.800 13.700 ;
        RECT 108.400 13.600 109.200 13.700 ;
        RECT 150.000 14.300 150.800 14.400 ;
        RECT 159.600 14.300 160.400 14.400 ;
        RECT 150.000 13.700 160.400 14.300 ;
        RECT 150.000 13.600 150.800 13.700 ;
        RECT 159.600 13.600 160.400 13.700 ;
        RECT 169.200 14.300 170.000 14.400 ;
        RECT 175.600 14.300 176.400 14.400 ;
        RECT 169.200 13.700 176.400 14.300 ;
        RECT 169.200 13.600 170.000 13.700 ;
        RECT 175.600 13.600 176.400 13.700 ;
        RECT 178.800 14.300 179.600 14.400 ;
        RECT 185.200 14.300 186.000 14.400 ;
        RECT 191.600 14.300 192.400 14.400 ;
        RECT 178.800 13.700 192.400 14.300 ;
        RECT 178.800 13.600 179.600 13.700 ;
        RECT 185.200 13.600 186.000 13.700 ;
        RECT 191.600 13.600 192.400 13.700 ;
        RECT 18.800 12.300 19.600 12.400 ;
        RECT 25.200 12.300 26.000 12.400 ;
        RECT 18.800 11.700 26.000 12.300 ;
        RECT 18.800 11.600 19.600 11.700 ;
        RECT 25.200 11.600 26.000 11.700 ;
        RECT 28.400 12.300 29.200 12.400 ;
        RECT 31.600 12.300 32.400 12.400 ;
        RECT 38.000 12.300 38.800 12.400 ;
        RECT 28.400 11.700 38.800 12.300 ;
        RECT 28.400 11.600 29.200 11.700 ;
        RECT 31.600 11.600 32.400 11.700 ;
        RECT 38.000 11.600 38.800 11.700 ;
        RECT 52.400 12.300 53.200 12.400 ;
        RECT 58.800 12.300 59.600 12.400 ;
        RECT 52.400 11.700 59.600 12.300 ;
        RECT 52.400 11.600 53.200 11.700 ;
        RECT 58.800 11.600 59.600 11.700 ;
        RECT 63.600 12.300 64.400 12.400 ;
        RECT 76.400 12.300 77.200 12.400 ;
        RECT 63.600 11.700 77.200 12.300 ;
        RECT 63.600 11.600 64.400 11.700 ;
        RECT 76.400 11.600 77.200 11.700 ;
        RECT 81.200 12.300 82.000 12.400 ;
        RECT 87.600 12.300 88.400 12.400 ;
        RECT 81.200 11.700 88.400 12.300 ;
        RECT 81.200 11.600 82.000 11.700 ;
        RECT 87.600 11.600 88.400 11.700 ;
        RECT 110.000 12.300 110.800 12.400 ;
        RECT 116.400 12.300 117.200 12.400 ;
        RECT 110.000 11.700 117.200 12.300 ;
        RECT 110.000 11.600 110.800 11.700 ;
        RECT 116.400 11.600 117.200 11.700 ;
        RECT 119.600 12.300 120.400 12.400 ;
        RECT 122.800 12.300 123.600 12.400 ;
        RECT 150.000 12.300 150.800 12.400 ;
        RECT 119.600 11.700 150.800 12.300 ;
        RECT 119.600 11.600 120.400 11.700 ;
        RECT 122.800 11.600 123.600 11.700 ;
        RECT 150.000 11.600 150.800 11.700 ;
        RECT 161.200 12.300 162.000 12.400 ;
        RECT 167.600 12.300 168.400 12.400 ;
        RECT 161.200 11.700 168.400 12.300 ;
        RECT 161.200 11.600 162.000 11.700 ;
        RECT 167.600 11.600 168.400 11.700 ;
        RECT 172.400 12.300 173.200 12.400 ;
        RECT 183.600 12.300 184.400 12.400 ;
        RECT 172.400 11.700 184.400 12.300 ;
        RECT 172.400 11.600 173.200 11.700 ;
        RECT 183.600 11.600 184.400 11.700 ;
        RECT 105.200 10.300 106.000 10.400 ;
        RECT 126.000 10.300 126.800 10.400 ;
        RECT 105.200 9.700 126.800 10.300 ;
        RECT 105.200 9.600 106.000 9.700 ;
        RECT 126.000 9.600 126.800 9.700 ;
      LAYER metal4 ;
        RECT 97.000 123.400 98.200 172.600 ;
        RECT 141.800 137.400 143.000 150.600 ;
        RECT 125.800 103.400 127.000 112.600 ;
        RECT 20.200 35.400 21.400 72.600 ;
        RECT 84.200 13.400 85.400 98.600 ;
        RECT 103.400 15.400 104.600 32.600 ;
        RECT 122.600 11.400 123.800 46.600 ;
  END
END address_gen
END LIBRARY

