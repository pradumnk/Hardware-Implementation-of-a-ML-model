magic
tech scmos
magscale 1 2
timestamp 1651681474
<< metal1 >>
rect 1352 1806 1358 1814
rect 1366 1806 1372 1814
rect 1380 1806 1386 1814
rect 1394 1806 1400 1814
rect 1869 1737 1884 1743
rect 573 1637 588 1643
rect 520 1606 526 1614
rect 534 1606 540 1614
rect 548 1606 554 1614
rect 562 1606 568 1614
rect 941 1517 956 1523
rect 1596 1506 1604 1516
rect 1380 1497 1395 1503
rect 1485 1497 1523 1503
rect 1533 1497 1548 1503
rect 1668 1497 1683 1503
rect 477 1477 515 1483
rect 596 1477 611 1483
rect 669 1477 684 1483
rect 788 1477 803 1483
rect 797 1457 803 1477
rect 868 1477 915 1483
rect 948 1477 963 1483
rect 1277 1477 1292 1483
rect 1309 1477 1388 1483
rect 1421 1477 1436 1483
rect 1740 1477 1764 1483
rect 1213 1457 1235 1463
rect 1352 1406 1358 1414
rect 1366 1406 1372 1414
rect 1380 1406 1386 1414
rect 1394 1406 1400 1414
rect 650 1376 652 1384
rect 781 1357 812 1363
rect 1668 1357 1699 1363
rect 1052 1344 1060 1348
rect 164 1337 179 1343
rect 356 1337 403 1343
rect 733 1337 748 1343
rect 1485 1337 1532 1343
rect 1572 1337 1587 1343
rect 621 1317 636 1323
rect 740 1317 755 1323
rect 765 1317 796 1323
rect 1236 1317 1251 1323
rect 1821 1317 1836 1323
rect 1316 1277 1331 1283
rect 458 1256 460 1264
rect 520 1206 526 1214
rect 534 1206 540 1214
rect 548 1206 554 1214
rect 562 1206 568 1214
rect 372 1176 374 1184
rect 420 1176 422 1184
rect 1658 1176 1660 1184
rect 996 1137 1011 1143
rect 1382 1136 1388 1144
rect 621 1117 636 1123
rect 685 1117 700 1123
rect 1476 1117 1491 1123
rect 1597 1117 1619 1123
rect 381 1097 412 1103
rect 717 1097 732 1103
rect 957 1097 979 1103
rect 1517 1097 1564 1103
rect 1581 1097 1596 1103
rect 964 1077 979 1083
rect 1533 1077 1548 1083
rect 1764 1077 1795 1083
rect 333 1057 348 1063
rect 1444 1057 1491 1063
rect 1629 1057 1644 1063
rect 1421 1037 1452 1043
rect 1352 1006 1358 1014
rect 1366 1006 1372 1014
rect 1380 1006 1386 1014
rect 1394 1006 1400 1014
rect 468 976 470 984
rect 1698 977 1740 983
rect 1917 977 1932 983
rect 92 957 124 963
rect 92 948 100 957
rect 349 957 387 963
rect 829 957 844 963
rect 1613 957 1651 963
rect 324 937 339 943
rect 429 937 451 943
rect 708 937 723 943
rect 1133 937 1148 943
rect 1357 937 1420 943
rect 45 917 68 923
rect 60 914 68 917
rect 285 917 323 923
rect 429 917 444 923
rect 525 917 540 923
rect 669 917 707 923
rect 813 917 851 923
rect 861 917 876 923
rect 996 917 1011 923
rect 1652 917 1683 923
rect 1732 917 1763 923
rect 1308 912 1316 916
rect 1156 877 1171 883
rect 520 806 526 814
rect 534 806 540 814
rect 548 806 554 814
rect 562 806 568 814
rect 925 737 948 743
rect 1245 737 1260 743
rect 157 697 195 703
rect 1325 697 1388 703
rect 1037 677 1052 683
rect 1277 677 1299 683
rect 1485 677 1500 683
rect 196 657 211 663
rect 260 657 291 663
rect 365 657 380 663
rect 628 657 675 663
rect 1485 657 1491 677
rect 1352 606 1358 614
rect 1366 606 1372 614
rect 1380 606 1386 614
rect 1394 606 1400 614
rect 724 557 755 563
rect 884 556 892 564
rect 1588 557 1603 563
rect 1812 556 1820 564
rect 1085 537 1164 543
rect 1229 537 1276 543
rect 1789 537 1804 543
rect 45 517 68 523
rect 60 514 68 517
rect 740 517 771 523
rect 781 517 803 523
rect 1133 517 1164 523
rect 1700 517 1715 523
rect 1837 523 1843 536
rect 1837 517 1859 523
rect 1556 497 1571 503
rect 1796 497 1811 503
rect 1588 477 1603 483
rect 1300 436 1302 444
rect 520 406 526 414
rect 534 406 540 414
rect 548 406 554 414
rect 562 406 568 414
rect 749 317 771 323
rect 948 317 963 323
rect 260 297 291 303
rect 301 297 339 303
rect 532 297 611 303
rect 1213 297 1251 303
rect 1261 297 1324 303
rect 372 277 387 283
rect 397 277 412 283
rect 484 277 499 283
rect 509 277 588 283
rect 493 257 499 277
rect 621 277 636 283
rect 1021 283 1027 296
rect 1005 277 1027 283
rect 1085 277 1123 283
rect 1708 277 1732 283
rect 1564 263 1572 272
rect 1564 257 1596 263
rect 1352 206 1358 214
rect 1366 206 1372 214
rect 1380 206 1386 214
rect 1394 206 1400 214
rect 1178 176 1180 184
rect 429 157 444 163
rect 1661 137 1692 143
rect 429 117 451 123
rect 461 117 524 123
rect 1388 117 1459 123
rect 1388 114 1396 117
rect 520 6 526 14
rect 534 6 540 14
rect 548 6 554 14
rect 562 6 568 14
<< m2contact >>
rect 1358 1806 1366 1814
rect 1372 1806 1380 1814
rect 1386 1806 1394 1814
rect 380 1776 388 1784
rect 668 1776 676 1784
rect 716 1776 724 1784
rect 764 1776 772 1784
rect 972 1776 980 1784
rect 1020 1776 1028 1784
rect 1292 1776 1300 1784
rect 1340 1776 1348 1784
rect 1628 1776 1636 1784
rect 1820 1776 1828 1784
rect 1884 1756 1892 1764
rect 12 1736 20 1744
rect 268 1736 276 1744
rect 412 1736 420 1744
rect 940 1736 948 1744
rect 1660 1736 1668 1744
rect 1884 1736 1892 1744
rect 284 1718 292 1726
rect 348 1716 356 1724
rect 460 1716 468 1724
rect 636 1716 644 1724
rect 684 1716 692 1724
rect 732 1716 740 1724
rect 908 1718 916 1726
rect 1004 1716 1012 1724
rect 1052 1716 1060 1724
rect 1132 1716 1140 1724
rect 1196 1718 1204 1726
rect 1260 1716 1268 1724
rect 1308 1716 1316 1724
rect 1468 1716 1476 1724
rect 1532 1718 1540 1726
rect 1596 1716 1604 1724
rect 1708 1716 1716 1724
rect 1836 1716 1844 1724
rect 1900 1716 1908 1724
rect 1404 1676 1412 1684
rect 1932 1676 1940 1684
rect 124 1636 132 1644
rect 156 1636 164 1644
rect 588 1636 596 1644
rect 780 1636 788 1644
rect 1068 1636 1076 1644
rect 526 1606 534 1614
rect 540 1606 548 1614
rect 554 1606 562 1614
rect 396 1576 404 1584
rect 1004 1576 1012 1584
rect 1132 1576 1140 1584
rect 1564 1536 1572 1544
rect 636 1516 644 1524
rect 748 1516 756 1524
rect 956 1516 964 1524
rect 1228 1516 1236 1524
rect 1324 1516 1332 1524
rect 1500 1516 1508 1524
rect 1596 1516 1604 1524
rect 140 1494 148 1502
rect 268 1496 276 1504
rect 332 1494 340 1502
rect 492 1496 500 1504
rect 524 1496 532 1504
rect 700 1496 708 1504
rect 732 1496 740 1504
rect 828 1496 836 1504
rect 892 1496 900 1504
rect 972 1496 980 1504
rect 1164 1496 1172 1504
rect 1196 1496 1204 1504
rect 1260 1496 1268 1504
rect 1372 1496 1380 1504
rect 1468 1496 1476 1504
rect 1548 1496 1556 1504
rect 1628 1496 1636 1504
rect 1660 1496 1668 1504
rect 1804 1494 1812 1502
rect 124 1476 132 1484
rect 172 1476 180 1484
rect 428 1480 436 1488
rect 444 1476 452 1484
rect 588 1476 596 1484
rect 684 1476 692 1484
rect 716 1476 724 1484
rect 780 1476 788 1484
rect 460 1456 468 1464
rect 540 1456 548 1464
rect 652 1456 660 1464
rect 684 1456 692 1464
rect 812 1476 820 1484
rect 860 1476 868 1484
rect 940 1476 948 1484
rect 1020 1476 1028 1484
rect 1180 1476 1188 1484
rect 1292 1476 1300 1484
rect 1388 1476 1396 1484
rect 1404 1476 1412 1484
rect 1436 1476 1444 1484
rect 1452 1476 1460 1484
rect 876 1456 884 1464
rect 940 1456 948 1464
rect 1436 1456 1444 1464
rect 1548 1456 1556 1464
rect 12 1436 20 1444
rect 204 1436 212 1444
rect 636 1436 644 1444
rect 748 1436 756 1444
rect 1932 1436 1940 1444
rect 1358 1406 1366 1414
rect 1372 1406 1380 1414
rect 1386 1406 1394 1414
rect 140 1376 148 1384
rect 316 1376 324 1384
rect 412 1376 420 1384
rect 652 1376 660 1384
rect 684 1376 692 1384
rect 844 1376 852 1384
rect 1036 1376 1044 1384
rect 1548 1376 1556 1384
rect 1708 1376 1716 1384
rect 156 1356 164 1364
rect 236 1356 244 1364
rect 252 1356 260 1364
rect 364 1356 372 1364
rect 428 1356 436 1364
rect 476 1356 484 1364
rect 508 1356 516 1364
rect 620 1356 628 1364
rect 1228 1356 1236 1364
rect 1324 1356 1332 1364
rect 1436 1356 1444 1364
rect 1452 1356 1460 1364
rect 1468 1356 1476 1364
rect 1564 1356 1572 1364
rect 60 1336 68 1344
rect 124 1336 132 1344
rect 156 1336 164 1344
rect 204 1336 212 1344
rect 268 1336 276 1344
rect 284 1336 292 1344
rect 348 1336 356 1344
rect 588 1336 596 1344
rect 668 1336 676 1344
rect 748 1336 756 1344
rect 828 1336 836 1344
rect 1004 1336 1012 1344
rect 1052 1336 1060 1344
rect 1308 1336 1316 1344
rect 1356 1336 1364 1344
rect 1532 1336 1540 1344
rect 1564 1336 1572 1344
rect 1612 1336 1620 1344
rect 1644 1336 1652 1344
rect 1724 1336 1732 1344
rect 1772 1336 1780 1344
rect 44 1316 52 1324
rect 92 1316 100 1324
rect 108 1316 116 1324
rect 188 1316 196 1324
rect 380 1316 388 1324
rect 444 1316 452 1324
rect 572 1316 580 1324
rect 636 1316 644 1324
rect 716 1316 724 1324
rect 732 1316 740 1324
rect 796 1316 804 1324
rect 956 1316 964 1324
rect 1100 1316 1108 1324
rect 1148 1316 1156 1324
rect 1228 1316 1236 1324
rect 1260 1316 1268 1324
rect 1372 1316 1380 1324
rect 1500 1316 1508 1324
rect 1516 1316 1524 1324
rect 1596 1316 1604 1324
rect 1740 1316 1748 1324
rect 1836 1316 1844 1324
rect 220 1296 228 1304
rect 300 1296 308 1304
rect 636 1296 644 1304
rect 684 1296 692 1304
rect 796 1296 804 1304
rect 1276 1296 1284 1304
rect 1628 1296 1636 1304
rect 1676 1296 1684 1304
rect 12 1276 20 1284
rect 1308 1276 1316 1284
rect 460 1256 468 1264
rect 492 1236 500 1244
rect 1292 1236 1300 1244
rect 1932 1236 1940 1244
rect 526 1206 534 1214
rect 540 1206 548 1214
rect 554 1206 562 1214
rect 364 1176 372 1184
rect 412 1176 420 1184
rect 460 1176 468 1184
rect 604 1176 612 1184
rect 1660 1176 1668 1184
rect 1852 1176 1860 1184
rect 1708 1156 1716 1164
rect 60 1136 68 1144
rect 476 1136 484 1144
rect 588 1136 596 1144
rect 988 1136 996 1144
rect 1388 1136 1396 1144
rect 1724 1136 1732 1144
rect 252 1116 260 1124
rect 444 1116 452 1124
rect 508 1116 516 1124
rect 636 1116 644 1124
rect 700 1116 708 1124
rect 732 1116 740 1124
rect 828 1116 836 1124
rect 844 1116 852 1124
rect 1468 1116 1476 1124
rect 1692 1116 1700 1124
rect 44 1096 52 1104
rect 188 1094 196 1102
rect 284 1096 292 1104
rect 412 1096 420 1104
rect 492 1096 500 1104
rect 604 1096 612 1104
rect 652 1096 660 1104
rect 732 1096 740 1104
rect 780 1096 788 1104
rect 876 1096 884 1104
rect 924 1096 932 1104
rect 1116 1096 1124 1104
rect 1196 1096 1204 1104
rect 1292 1094 1300 1102
rect 1564 1096 1572 1104
rect 1596 1096 1604 1104
rect 1644 1096 1652 1104
rect 1708 1096 1716 1104
rect 1804 1096 1812 1104
rect 1884 1096 1892 1104
rect 12 1076 20 1084
rect 172 1076 180 1084
rect 300 1076 308 1084
rect 396 1076 404 1084
rect 636 1076 644 1084
rect 700 1076 708 1084
rect 796 1076 804 1084
rect 860 1076 868 1084
rect 892 1076 900 1084
rect 940 1076 948 1084
rect 956 1076 964 1084
rect 1100 1076 1108 1084
rect 1260 1076 1268 1084
rect 1548 1076 1556 1084
rect 1756 1076 1764 1084
rect 1916 1076 1924 1084
rect 316 1056 324 1064
rect 348 1056 356 1064
rect 748 1056 756 1064
rect 908 1056 916 1064
rect 988 1056 996 1064
rect 1228 1056 1236 1064
rect 1436 1056 1444 1064
rect 1644 1056 1652 1064
rect 1676 1056 1684 1064
rect 1772 1056 1780 1064
rect 764 1036 772 1044
rect 828 1036 836 1044
rect 1212 1036 1220 1044
rect 1452 1036 1460 1044
rect 1358 1006 1366 1014
rect 1372 1006 1380 1014
rect 1386 1006 1394 1014
rect 380 976 388 984
rect 460 976 468 984
rect 492 976 500 984
rect 636 976 644 984
rect 748 976 756 984
rect 892 976 900 984
rect 1116 976 1124 984
rect 1228 976 1236 984
rect 1740 976 1748 984
rect 1932 976 1940 984
rect 124 956 132 964
rect 396 956 404 964
rect 412 956 420 964
rect 732 956 740 964
rect 844 956 852 964
rect 876 956 884 964
rect 1148 956 1156 964
rect 1180 956 1188 964
rect 1244 956 1252 964
rect 1372 956 1380 964
rect 1436 956 1444 964
rect 1532 956 1540 964
rect 1596 956 1604 964
rect 1820 956 1828 964
rect 172 936 180 944
rect 252 936 260 944
rect 316 936 324 944
rect 588 936 596 944
rect 652 936 660 944
rect 700 936 708 944
rect 1148 936 1156 944
rect 1212 936 1220 944
rect 1340 936 1348 944
rect 1420 936 1428 944
rect 1452 936 1460 944
rect 1484 936 1492 944
rect 1516 936 1524 944
rect 1564 936 1572 944
rect 1660 936 1668 944
rect 1788 936 1796 944
rect 188 918 196 926
rect 268 916 276 924
rect 364 916 372 924
rect 444 916 452 924
rect 540 916 548 924
rect 604 916 612 924
rect 780 916 788 924
rect 796 916 804 924
rect 876 916 884 924
rect 956 916 964 924
rect 988 916 996 924
rect 1084 916 1092 924
rect 1196 916 1204 924
rect 1260 916 1268 924
rect 1292 916 1300 924
rect 1308 916 1316 924
rect 1324 916 1332 924
rect 1500 916 1508 924
rect 1580 916 1588 924
rect 1644 916 1652 924
rect 1724 916 1732 924
rect 1836 916 1844 924
rect 1884 916 1892 924
rect 300 896 308 904
rect 476 896 484 904
rect 684 896 692 904
rect 1468 896 1476 904
rect 12 876 20 884
rect 1148 876 1156 884
rect 1276 876 1284 884
rect 1868 876 1876 884
rect 60 836 68 844
rect 1532 836 1540 844
rect 1804 836 1812 844
rect 526 806 534 814
rect 540 806 548 814
rect 554 806 562 814
rect 92 776 100 784
rect 300 776 308 784
rect 684 776 692 784
rect 860 776 868 784
rect 1916 776 1924 784
rect 76 736 84 744
rect 604 736 612 744
rect 1260 736 1268 744
rect 108 716 116 724
rect 172 716 180 724
rect 268 716 276 724
rect 364 716 372 724
rect 396 716 404 724
rect 940 716 948 724
rect 1340 716 1348 724
rect 1468 716 1476 724
rect 1532 716 1540 724
rect 44 696 52 704
rect 92 696 100 704
rect 140 696 148 704
rect 332 696 340 704
rect 380 696 388 704
rect 476 694 484 702
rect 732 696 740 704
rect 892 696 900 704
rect 972 696 980 704
rect 1052 696 1060 704
rect 1116 694 1124 702
rect 1276 696 1284 704
rect 1308 696 1316 704
rect 1388 696 1396 704
rect 1420 696 1428 704
rect 1452 696 1460 704
rect 1660 696 1668 704
rect 1788 694 1796 702
rect 12 676 20 684
rect 124 676 132 684
rect 236 676 244 684
rect 300 676 308 684
rect 316 676 324 684
rect 748 676 756 684
rect 956 676 964 684
rect 988 676 996 684
rect 1020 676 1028 684
rect 1052 676 1060 684
rect 1084 676 1092 684
rect 1404 676 1412 684
rect 188 656 196 664
rect 220 656 228 664
rect 380 656 388 664
rect 412 656 420 664
rect 476 656 484 664
rect 620 656 628 664
rect 1004 656 1012 664
rect 1260 656 1268 664
rect 1500 676 1508 684
rect 1756 676 1764 684
rect 1676 656 1684 664
rect 700 636 708 644
rect 1532 636 1540 644
rect 1548 636 1556 644
rect 1358 606 1366 614
rect 1372 606 1380 614
rect 1386 606 1394 614
rect 60 576 68 584
rect 300 576 308 584
rect 1052 576 1060 584
rect 1228 576 1236 584
rect 1388 576 1396 584
rect 1452 576 1460 584
rect 1644 576 1652 584
rect 1740 576 1748 584
rect 796 556 804 564
rect 892 556 900 564
rect 1100 556 1108 564
rect 1228 556 1236 564
rect 1580 556 1588 564
rect 1692 556 1700 564
rect 1804 556 1812 564
rect 172 536 180 544
rect 220 536 228 544
rect 252 536 260 544
rect 268 532 276 540
rect 316 536 324 544
rect 444 536 452 544
rect 524 536 532 544
rect 700 536 708 544
rect 828 536 836 544
rect 860 536 868 544
rect 908 536 916 544
rect 1164 536 1172 544
rect 1276 536 1284 544
rect 1436 536 1444 544
rect 1484 536 1492 544
rect 1500 536 1508 544
rect 1804 536 1812 544
rect 1836 536 1844 544
rect 1884 536 1892 544
rect 188 518 196 526
rect 572 516 580 524
rect 732 516 740 524
rect 844 516 852 524
rect 1164 516 1172 524
rect 1212 516 1220 524
rect 1292 516 1300 524
rect 1420 516 1428 524
rect 1516 516 1524 524
rect 1580 516 1588 524
rect 1660 516 1668 524
rect 1692 516 1700 524
rect 1724 516 1732 524
rect 1772 516 1780 524
rect 1900 516 1908 524
rect 732 496 740 504
rect 892 496 900 504
rect 1052 496 1060 504
rect 1324 496 1332 504
rect 1452 496 1460 504
rect 1548 496 1556 504
rect 1676 496 1684 504
rect 1788 496 1796 504
rect 12 476 20 484
rect 1580 476 1588 484
rect 1644 476 1652 484
rect 1932 476 1940 484
rect 684 436 692 444
rect 1020 436 1028 444
rect 1292 436 1300 444
rect 1612 436 1620 444
rect 526 406 534 414
rect 540 406 548 414
rect 554 406 562 414
rect 732 376 740 384
rect 1532 376 1540 384
rect 1900 376 1908 384
rect 684 336 692 344
rect 716 336 724 344
rect 204 316 212 324
rect 316 316 324 324
rect 412 316 420 324
rect 428 316 436 324
rect 588 316 596 324
rect 940 316 948 324
rect 1164 316 1172 324
rect 1228 316 1236 324
rect 140 294 148 302
rect 236 296 244 304
rect 252 296 260 304
rect 348 296 356 304
rect 460 296 468 304
rect 524 296 532 304
rect 652 296 660 304
rect 732 296 740 304
rect 796 296 804 304
rect 828 296 836 304
rect 908 296 916 304
rect 988 296 996 304
rect 1020 296 1028 304
rect 1084 296 1092 304
rect 1132 296 1140 304
rect 1196 296 1204 304
rect 1324 296 1332 304
rect 172 276 180 284
rect 252 276 260 284
rect 364 276 372 284
rect 412 276 420 284
rect 476 276 484 284
rect 268 256 276 264
rect 588 276 596 284
rect 636 276 644 284
rect 812 276 820 284
rect 844 276 852 284
rect 892 276 900 284
rect 924 276 932 284
rect 972 276 980 284
rect 1388 294 1396 302
rect 1596 296 1604 304
rect 1660 294 1668 302
rect 1788 296 1796 304
rect 1036 276 1044 284
rect 1164 276 1172 284
rect 1180 276 1188 284
rect 1420 276 1428 284
rect 876 256 884 264
rect 1068 256 1076 264
rect 1100 256 1108 264
rect 1276 256 1284 264
rect 1596 256 1604 264
rect 12 236 20 244
rect 204 236 212 244
rect 428 236 436 244
rect 860 236 868 244
rect 1052 236 1060 244
rect 1516 236 1524 244
rect 1358 206 1366 214
rect 1372 206 1380 214
rect 1386 206 1394 214
rect 60 176 68 184
rect 716 176 724 184
rect 972 176 980 184
rect 1180 176 1188 184
rect 1388 176 1396 184
rect 1804 176 1812 184
rect 1884 176 1892 184
rect 252 156 260 164
rect 444 156 452 164
rect 476 156 484 164
rect 1644 156 1652 164
rect 1724 156 1732 164
rect 1740 156 1748 164
rect 1868 156 1876 164
rect 172 136 180 144
rect 284 136 292 144
rect 348 132 356 140
rect 364 136 372 144
rect 396 136 404 144
rect 556 136 564 144
rect 1068 136 1076 144
rect 1196 136 1204 144
rect 1228 136 1236 144
rect 1692 136 1700 144
rect 1756 136 1764 144
rect 1788 136 1796 144
rect 1852 136 1860 144
rect 1900 136 1908 144
rect 44 116 52 124
rect 188 118 196 126
rect 252 116 260 124
rect 300 116 308 124
rect 316 116 324 124
rect 380 116 388 124
rect 524 116 532 124
rect 588 118 596 126
rect 764 116 772 124
rect 780 116 788 124
rect 828 116 836 124
rect 876 116 884 124
rect 924 116 932 124
rect 1084 116 1092 124
rect 1260 118 1268 126
rect 1500 116 1508 124
rect 1548 116 1556 124
rect 1596 116 1604 124
rect 1676 116 1684 124
rect 1724 116 1732 124
rect 1836 116 1844 124
rect 1916 116 1924 124
rect 1164 96 1172 104
rect 12 76 20 84
rect 732 36 740 44
rect 812 36 820 44
rect 860 36 868 44
rect 908 36 916 44
rect 956 36 964 44
rect 1484 36 1492 44
rect 1532 36 1540 44
rect 1580 36 1588 44
rect 1628 36 1636 44
rect 526 6 534 14
rect 540 6 548 14
rect 554 6 562 14
<< metal2 >>
rect 365 1837 387 1843
rect 381 1784 387 1837
rect 637 1804 643 1843
rect 685 1804 691 1843
rect 749 1837 771 1843
rect 669 1784 675 1796
rect 717 1784 723 1796
rect 765 1784 771 1837
rect 973 1837 995 1843
rect 1021 1837 1043 1843
rect 1277 1837 1299 1843
rect 973 1784 979 1837
rect 1021 1784 1027 1837
rect 1293 1784 1299 1837
rect 1325 1783 1331 1843
rect 1613 1837 1635 1843
rect 1352 1806 1358 1814
rect 1366 1806 1372 1814
rect 1380 1806 1386 1814
rect 1394 1806 1400 1814
rect 1629 1784 1635 1837
rect 1325 1777 1340 1783
rect 1821 1744 1827 1776
rect 1853 1764 1859 1843
rect 13 1704 19 1736
rect 125 1504 131 1636
rect 157 1604 163 1636
rect 125 1484 131 1496
rect 13 1324 19 1436
rect 93 1324 99 1436
rect 141 1384 147 1494
rect 125 1304 131 1336
rect 157 1324 163 1336
rect 13 1284 19 1296
rect 61 1104 67 1136
rect 13 1084 19 1096
rect 173 1084 179 1476
rect 237 1364 243 1596
rect 269 1504 275 1736
rect 285 1664 291 1718
rect 1133 1724 1139 1736
rect 349 1604 355 1716
rect 461 1664 467 1716
rect 397 1584 403 1656
rect 520 1606 526 1614
rect 534 1606 540 1614
rect 548 1606 554 1614
rect 562 1606 568 1614
rect 589 1524 595 1636
rect 637 1524 643 1716
rect 685 1524 691 1716
rect 733 1664 739 1716
rect 909 1704 915 1718
rect 1469 1724 1475 1736
rect 621 1517 636 1523
rect 413 1480 428 1483
rect 413 1477 435 1480
rect 205 1344 211 1356
rect 237 1344 243 1356
rect 189 1304 195 1316
rect 301 1304 307 1436
rect 317 1384 323 1456
rect 413 1384 419 1477
rect 445 1464 451 1476
rect 493 1464 499 1496
rect 461 1444 467 1456
rect 541 1444 547 1456
rect 372 1357 387 1363
rect 349 1344 355 1356
rect 381 1324 387 1357
rect 189 1102 195 1116
rect 221 1084 227 1296
rect 365 1284 371 1296
rect 365 1184 371 1276
rect 381 1244 387 1316
rect 429 1164 435 1356
rect 589 1344 595 1476
rect 621 1384 627 1517
rect 653 1464 659 1516
rect 701 1504 707 1656
rect 781 1644 787 1656
rect 781 1484 787 1636
rect 1005 1584 1011 1696
rect 877 1497 892 1503
rect 877 1464 883 1497
rect 957 1503 963 1516
rect 957 1497 972 1503
rect 941 1484 947 1496
rect 1021 1484 1027 1676
rect 1021 1464 1027 1476
rect 621 1364 627 1376
rect 637 1364 643 1436
rect 653 1384 659 1436
rect 685 1384 691 1456
rect 749 1344 755 1436
rect 836 1337 851 1343
rect 445 1324 451 1336
rect 589 1324 595 1336
rect 573 1284 579 1316
rect 669 1303 675 1336
rect 669 1297 684 1303
rect 637 1284 643 1296
rect 717 1284 723 1316
rect 461 1184 467 1236
rect 173 944 179 1076
rect 285 1004 291 1056
rect 253 944 259 956
rect 189 926 195 936
rect 13 884 19 896
rect 68 837 83 843
rect 77 744 83 837
rect 93 784 99 916
rect 269 824 275 916
rect 141 704 147 716
rect 13 684 19 696
rect 125 564 131 676
rect 141 584 147 696
rect 237 684 243 696
rect 269 664 275 716
rect 13 484 19 496
rect 173 284 179 536
rect 189 526 195 656
rect 253 544 259 556
rect 269 540 275 576
rect 285 564 291 996
rect 301 904 307 1076
rect 381 984 387 1136
rect 397 1064 403 1076
rect 397 964 403 1056
rect 413 984 419 1096
rect 445 1084 451 1116
rect 413 924 419 956
rect 477 904 483 1116
rect 493 1104 499 1236
rect 520 1206 526 1214
rect 534 1206 540 1214
rect 548 1206 554 1214
rect 562 1206 568 1214
rect 605 1184 611 1276
rect 493 984 499 1076
rect 541 904 547 916
rect 301 844 307 896
rect 301 784 307 816
rect 365 724 371 836
rect 520 806 526 814
rect 534 806 540 814
rect 548 806 554 814
rect 562 806 568 814
rect 477 702 483 716
rect 605 704 611 736
rect 317 684 323 696
rect 333 664 339 696
rect 381 684 387 696
rect 621 664 627 1156
rect 637 1084 643 1116
rect 653 1104 659 1256
rect 637 1024 643 1076
rect 637 964 643 976
rect 653 944 659 996
rect 685 904 691 976
rect 701 964 707 1076
rect 749 1064 755 1336
rect 845 1304 851 1337
rect 781 1104 787 1276
rect 797 1244 803 1296
rect 845 1124 851 1296
rect 877 1284 883 1456
rect 941 1164 947 1456
rect 829 1104 835 1116
rect 733 1057 748 1063
rect 733 964 739 1057
rect 797 1044 803 1076
rect 845 1044 851 1116
rect 925 1104 931 1116
rect 941 1084 947 1096
rect 861 1064 867 1076
rect 973 1044 979 1456
rect 1037 1304 1043 1376
rect 1053 1344 1059 1716
rect 1069 1484 1075 1636
rect 1133 1584 1139 1716
rect 1197 1504 1203 1718
rect 1261 1604 1267 1716
rect 1309 1684 1315 1716
rect 1165 1484 1171 1496
rect 1181 1484 1187 1496
rect 1293 1484 1299 1596
rect 1181 1463 1187 1476
rect 1165 1457 1187 1463
rect 1101 1324 1107 1336
rect 989 1144 995 1236
rect 989 1064 995 1136
rect 1101 1104 1107 1316
rect 1165 1144 1171 1457
rect 1197 1184 1203 1356
rect 1309 1344 1315 1676
rect 1325 1464 1331 1516
rect 1373 1444 1379 1496
rect 1389 1484 1395 1496
rect 1453 1484 1459 1496
rect 1469 1463 1475 1496
rect 1453 1457 1475 1463
rect 1352 1406 1358 1414
rect 1366 1406 1372 1414
rect 1380 1406 1386 1414
rect 1394 1406 1400 1414
rect 1437 1364 1443 1436
rect 1453 1364 1459 1457
rect 1533 1443 1539 1718
rect 1549 1464 1555 1476
rect 1565 1464 1571 1536
rect 1597 1524 1603 1716
rect 1629 1504 1635 1736
rect 1533 1437 1555 1443
rect 1549 1384 1555 1437
rect 1469 1364 1475 1376
rect 1309 1324 1315 1336
rect 1261 1284 1267 1316
rect 1325 1304 1331 1356
rect 1357 1324 1363 1336
rect 1373 1324 1379 1336
rect 1117 1104 1123 1116
rect 1197 1104 1203 1136
rect 1101 1084 1107 1096
rect 749 984 755 1036
rect 765 924 771 1036
rect 829 964 835 1036
rect 845 964 851 976
rect 781 904 787 916
rect 733 784 739 896
rect 861 784 867 816
rect 733 704 739 776
rect 893 704 899 896
rect 301 584 307 656
rect 445 544 451 556
rect 477 544 483 656
rect 701 544 707 636
rect 749 564 755 676
rect 804 557 819 563
rect 749 544 755 556
rect 205 324 211 356
rect 253 324 259 536
rect 520 406 526 414
rect 534 406 540 414
rect 548 406 554 414
rect 562 406 568 414
rect 701 364 707 536
rect 813 524 819 557
rect 909 544 915 1036
rect 957 824 963 916
rect 1085 904 1091 916
rect 1101 823 1107 1076
rect 1117 984 1123 1076
rect 1229 1064 1235 1176
rect 1293 1144 1299 1236
rect 1389 1144 1395 1276
rect 1469 1184 1475 1356
rect 1501 1324 1507 1356
rect 1613 1344 1619 1356
rect 1645 1344 1651 1516
rect 1725 1423 1731 1496
rect 1709 1417 1731 1423
rect 1709 1384 1715 1417
rect 1565 1324 1571 1336
rect 1597 1324 1603 1336
rect 1645 1303 1651 1336
rect 1636 1297 1651 1303
rect 1293 1102 1299 1116
rect 1261 1084 1267 1096
rect 1469 1084 1475 1116
rect 1549 1084 1555 1116
rect 1597 1104 1603 1296
rect 1213 1024 1219 1036
rect 1229 984 1235 1036
rect 1261 963 1267 1056
rect 1352 1006 1358 1014
rect 1366 1006 1372 1014
rect 1380 1006 1386 1014
rect 1394 1006 1400 1014
rect 1373 964 1379 976
rect 1252 957 1267 963
rect 1092 817 1107 823
rect 733 384 739 496
rect 813 444 819 516
rect 317 324 323 356
rect 429 324 435 356
rect 733 324 739 376
rect 349 304 355 316
rect 237 284 243 296
rect 45 124 51 236
rect 173 144 179 276
rect 253 264 259 276
rect 269 264 275 276
rect 205 204 211 236
rect 253 164 259 196
rect 269 123 275 256
rect 301 184 307 256
rect 301 164 307 176
rect 285 124 291 136
rect 301 124 307 156
rect 349 140 355 296
rect 365 244 371 276
rect 365 144 371 236
rect 269 117 284 123
rect 13 84 19 96
rect 349 -17 355 132
rect 381 124 387 256
rect 429 184 435 236
rect 445 164 451 316
rect 653 304 659 316
rect 477 164 483 176
rect 637 164 643 276
rect 717 184 723 316
rect 733 264 739 296
rect 813 284 819 436
rect 829 304 835 536
rect 861 524 867 536
rect 845 484 851 516
rect 941 504 947 716
rect 957 664 963 676
rect 973 644 979 696
rect 989 684 995 696
rect 1085 684 1091 816
rect 1117 684 1123 694
rect 1053 644 1059 676
rect 1053 584 1059 636
rect 845 284 851 476
rect 893 304 899 496
rect 941 324 947 496
rect 1053 484 1059 496
rect 1021 324 1027 436
rect 1149 323 1155 876
rect 1165 443 1171 516
rect 1181 464 1187 956
rect 1293 924 1299 936
rect 1373 924 1379 956
rect 1421 944 1427 1016
rect 1437 964 1443 996
rect 1453 964 1459 1036
rect 1437 944 1443 956
rect 1277 804 1283 876
rect 1325 804 1331 916
rect 1469 904 1475 1076
rect 1485 944 1491 956
rect 1565 944 1571 1096
rect 1629 1084 1635 1296
rect 1661 1184 1667 1336
rect 1741 1324 1747 1416
rect 1709 1124 1715 1156
rect 1645 1064 1651 1076
rect 1677 1064 1683 1116
rect 1693 984 1699 1116
rect 1709 1004 1715 1096
rect 1725 1044 1731 1136
rect 1741 1084 1747 1316
rect 1773 1284 1779 1336
rect 1773 1164 1779 1256
rect 1837 1243 1843 1316
rect 1853 1264 1859 1756
rect 1885 1723 1891 1736
rect 1885 1717 1900 1723
rect 1933 1684 1939 1696
rect 1933 1424 1939 1436
rect 1837 1237 1859 1243
rect 1853 1184 1859 1237
rect 1757 1063 1763 1076
rect 1773 1064 1779 1156
rect 1741 1057 1763 1063
rect 1597 964 1603 976
rect 1565 924 1571 936
rect 1581 924 1587 936
rect 1725 924 1731 1036
rect 1741 984 1747 1057
rect 1805 1024 1811 1096
rect 1885 1084 1891 1096
rect 1917 1084 1923 1096
rect 1933 1064 1939 1236
rect 1229 584 1235 796
rect 1533 744 1539 836
rect 1261 664 1267 736
rect 1517 717 1532 723
rect 1309 644 1315 696
rect 1412 677 1427 683
rect 1229 524 1235 556
rect 1277 544 1283 576
rect 1293 524 1299 636
rect 1352 606 1358 614
rect 1366 606 1372 614
rect 1380 606 1386 614
rect 1394 606 1400 614
rect 1389 564 1395 576
rect 1421 564 1427 677
rect 1501 644 1507 676
rect 1517 664 1523 717
rect 1437 544 1443 556
rect 1165 437 1187 443
rect 1149 317 1164 323
rect 989 304 995 316
rect 893 284 899 296
rect 909 284 915 296
rect 989 284 995 296
rect 1133 284 1139 296
rect 1181 284 1187 437
rect 1213 303 1219 516
rect 1421 504 1427 516
rect 1469 503 1475 576
rect 1501 544 1507 636
rect 1485 504 1491 536
rect 1460 497 1475 503
rect 1204 297 1219 303
rect 1229 284 1235 316
rect 397 144 403 156
rect 637 124 643 156
rect 717 144 723 176
rect 781 124 787 136
rect 813 124 819 276
rect 861 144 867 236
rect 893 184 899 276
rect 925 264 931 276
rect 973 264 979 276
rect 829 124 835 136
rect 925 124 931 176
rect 1053 104 1059 236
rect 1069 144 1075 156
rect 1085 124 1091 136
rect 1101 124 1107 256
rect 1181 184 1187 276
rect 1293 264 1299 436
rect 1421 284 1427 296
rect 1352 206 1358 214
rect 1366 206 1372 214
rect 1380 206 1386 214
rect 1394 206 1400 214
rect 1165 124 1171 176
rect 1421 164 1427 276
rect 1229 144 1235 156
rect 1501 144 1507 536
rect 1517 524 1523 656
rect 1533 604 1539 636
rect 1581 524 1587 536
rect 1517 284 1523 516
rect 1533 384 1539 516
rect 1597 304 1603 616
rect 1645 584 1651 916
rect 1821 903 1827 956
rect 1837 924 1843 996
rect 1885 984 1891 1056
rect 1885 924 1891 976
rect 1821 897 1843 903
rect 1789 702 1795 736
rect 1677 624 1683 656
rect 1757 624 1763 676
rect 1693 564 1699 596
rect 1805 583 1811 836
rect 1805 577 1827 583
rect 1661 524 1667 536
rect 1725 524 1731 556
rect 1693 503 1699 516
rect 1684 497 1699 503
rect 1773 503 1779 516
rect 1789 504 1795 516
rect 1773 497 1788 503
rect 1197 124 1203 136
rect 1165 104 1171 116
rect 1261 104 1267 118
rect 1517 123 1523 236
rect 1549 124 1555 276
rect 1597 164 1603 256
rect 1597 124 1603 136
rect 1613 124 1619 436
rect 1789 284 1795 296
rect 1725 164 1731 236
rect 1805 184 1811 296
rect 1821 164 1827 577
rect 1837 544 1843 897
rect 1869 884 1875 896
rect 1917 784 1923 996
rect 1837 384 1843 536
rect 1933 484 1939 496
rect 1869 164 1875 256
rect 1885 184 1891 276
rect 1677 124 1683 156
rect 1901 144 1907 156
rect 1917 124 1923 136
rect 1508 117 1523 123
rect 520 6 526 14
rect 534 6 540 14
rect 548 6 554 14
rect 562 6 568 14
rect 333 -23 355 -17
rect 733 -23 739 36
rect 813 -17 819 36
rect 861 -17 867 36
rect 909 -17 915 36
rect 957 -17 963 36
rect 1485 24 1491 36
rect 1533 24 1539 36
rect 1581 24 1587 36
rect 797 -23 819 -17
rect 845 -23 867 -17
rect 893 -23 915 -17
rect 941 -23 963 -17
rect 1453 -23 1459 16
rect 1501 -23 1507 16
rect 1549 -23 1555 16
rect 1629 -17 1635 36
rect 1613 -23 1635 -17
<< m3contact >>
rect 636 1796 644 1804
rect 668 1796 676 1804
rect 684 1796 692 1804
rect 716 1796 724 1804
rect 1358 1806 1366 1814
rect 1372 1806 1380 1814
rect 1386 1806 1394 1814
rect 1852 1756 1860 1764
rect 1884 1756 1892 1764
rect 268 1736 276 1744
rect 412 1736 420 1744
rect 940 1736 948 1744
rect 1132 1736 1140 1744
rect 1468 1736 1476 1744
rect 1628 1736 1636 1744
rect 1660 1736 1668 1744
rect 1820 1736 1828 1744
rect 12 1696 20 1704
rect 156 1596 164 1604
rect 236 1596 244 1604
rect 124 1496 132 1504
rect 92 1436 100 1444
rect 60 1336 68 1344
rect 156 1356 164 1364
rect 12 1316 20 1324
rect 44 1316 52 1324
rect 108 1316 116 1324
rect 156 1316 164 1324
rect 12 1296 20 1304
rect 124 1296 132 1304
rect 12 1096 20 1104
rect 44 1096 52 1104
rect 60 1096 68 1104
rect 204 1436 212 1444
rect 284 1656 292 1664
rect 396 1656 404 1664
rect 460 1656 468 1664
rect 348 1596 356 1604
rect 526 1606 534 1614
rect 540 1606 548 1614
rect 554 1606 562 1614
rect 1004 1716 1012 1724
rect 908 1696 916 1704
rect 1004 1696 1012 1704
rect 700 1656 708 1664
rect 732 1656 740 1664
rect 780 1656 788 1664
rect 588 1516 596 1524
rect 268 1496 276 1504
rect 332 1502 340 1504
rect 332 1496 340 1502
rect 524 1496 532 1504
rect 316 1456 324 1464
rect 300 1436 308 1444
rect 204 1356 212 1364
rect 252 1356 260 1364
rect 236 1336 244 1344
rect 268 1336 276 1344
rect 284 1336 292 1344
rect 444 1456 452 1464
rect 492 1456 500 1464
rect 460 1436 468 1444
rect 540 1436 548 1444
rect 348 1356 356 1364
rect 476 1356 484 1364
rect 508 1356 516 1364
rect 188 1296 196 1304
rect 364 1296 372 1304
rect 188 1116 196 1124
rect 364 1276 372 1284
rect 380 1236 388 1244
rect 412 1176 420 1184
rect 652 1516 660 1524
rect 684 1516 692 1524
rect 748 1516 756 1524
rect 732 1496 740 1504
rect 1020 1676 1028 1684
rect 828 1496 836 1504
rect 684 1476 692 1484
rect 716 1476 724 1484
rect 812 1476 820 1484
rect 860 1476 868 1484
rect 940 1496 948 1504
rect 972 1456 980 1464
rect 1020 1456 1028 1464
rect 652 1436 660 1444
rect 620 1376 628 1384
rect 636 1356 644 1364
rect 844 1376 852 1384
rect 444 1336 452 1344
rect 588 1316 596 1324
rect 636 1316 644 1324
rect 732 1316 740 1324
rect 684 1296 692 1304
rect 572 1276 580 1284
rect 604 1276 612 1284
rect 636 1276 644 1284
rect 716 1276 724 1284
rect 460 1256 468 1264
rect 460 1236 468 1244
rect 428 1156 436 1164
rect 380 1136 388 1144
rect 476 1136 484 1144
rect 252 1116 260 1124
rect 284 1096 292 1104
rect 220 1076 228 1084
rect 300 1076 308 1084
rect 124 956 132 964
rect 284 1056 292 1064
rect 284 996 292 1004
rect 252 956 260 964
rect 188 936 196 944
rect 92 916 100 924
rect 12 896 20 904
rect 268 816 276 824
rect 108 716 116 724
rect 140 716 148 724
rect 172 716 180 724
rect 12 696 20 704
rect 44 696 52 704
rect 92 696 100 704
rect 236 696 244 704
rect 60 576 68 584
rect 220 656 228 664
rect 268 656 276 664
rect 140 576 148 584
rect 124 556 132 564
rect 12 496 20 504
rect 140 302 148 304
rect 140 296 148 302
rect 268 576 276 584
rect 252 556 260 564
rect 220 536 228 544
rect 316 1056 324 1064
rect 348 1056 356 1064
rect 476 1116 484 1124
rect 396 1056 404 1064
rect 444 1076 452 1084
rect 412 976 420 984
rect 460 976 468 984
rect 316 936 324 944
rect 364 916 372 924
rect 412 916 420 924
rect 444 916 452 924
rect 526 1206 534 1214
rect 540 1206 548 1214
rect 554 1206 562 1214
rect 652 1256 660 1264
rect 620 1156 628 1164
rect 588 1136 596 1144
rect 508 1116 516 1124
rect 604 1096 612 1104
rect 492 1076 500 1084
rect 588 936 596 944
rect 604 916 612 924
rect 540 896 548 904
rect 300 836 308 844
rect 364 836 372 844
rect 300 816 308 824
rect 526 806 534 814
rect 540 806 548 814
rect 554 806 562 814
rect 396 716 404 724
rect 476 716 484 724
rect 316 696 324 704
rect 300 676 308 684
rect 604 696 612 704
rect 380 676 388 684
rect 636 1116 644 1124
rect 700 1116 708 1124
rect 732 1116 740 1124
rect 652 1096 660 1104
rect 732 1096 740 1104
rect 636 1016 644 1024
rect 652 996 660 1004
rect 636 956 644 964
rect 684 976 692 984
rect 796 1316 804 1324
rect 844 1296 852 1304
rect 780 1276 788 1284
rect 796 1236 804 1244
rect 876 1276 884 1284
rect 956 1316 964 1324
rect 940 1156 948 1164
rect 924 1116 932 1124
rect 828 1096 836 1104
rect 876 1096 884 1104
rect 940 1096 948 1104
rect 892 1076 900 1084
rect 956 1076 964 1084
rect 860 1056 868 1064
rect 908 1056 916 1064
rect 1004 1336 1012 1344
rect 1308 1676 1316 1684
rect 1404 1676 1412 1684
rect 1260 1596 1268 1604
rect 1292 1596 1300 1604
rect 1228 1516 1236 1524
rect 1180 1496 1188 1504
rect 1260 1496 1268 1504
rect 1068 1476 1076 1484
rect 1164 1476 1172 1484
rect 1292 1476 1300 1484
rect 1100 1336 1108 1344
rect 1148 1316 1156 1324
rect 1036 1296 1044 1304
rect 988 1236 996 1244
rect 1196 1356 1204 1364
rect 1228 1356 1236 1364
rect 1500 1516 1508 1524
rect 1372 1496 1380 1504
rect 1388 1496 1396 1504
rect 1452 1496 1460 1504
rect 1324 1456 1332 1464
rect 1404 1476 1412 1484
rect 1436 1476 1444 1484
rect 1436 1456 1444 1464
rect 1372 1436 1380 1444
rect 1436 1436 1444 1444
rect 1358 1406 1366 1414
rect 1372 1406 1380 1414
rect 1386 1406 1394 1414
rect 1548 1496 1556 1504
rect 1548 1476 1556 1484
rect 1708 1716 1716 1724
rect 1836 1716 1844 1724
rect 1644 1516 1652 1524
rect 1564 1456 1572 1464
rect 1468 1376 1476 1384
rect 1452 1356 1460 1364
rect 1500 1356 1508 1364
rect 1564 1356 1572 1364
rect 1612 1356 1620 1364
rect 1228 1316 1236 1324
rect 1308 1316 1316 1324
rect 1372 1336 1380 1344
rect 1356 1316 1364 1324
rect 1276 1296 1284 1304
rect 1324 1296 1332 1304
rect 1260 1276 1268 1284
rect 1308 1276 1316 1284
rect 1388 1276 1396 1284
rect 1196 1176 1204 1184
rect 1228 1176 1236 1184
rect 1164 1136 1172 1144
rect 1196 1136 1204 1144
rect 1116 1116 1124 1124
rect 1100 1096 1108 1104
rect 1116 1076 1124 1084
rect 748 1036 756 1044
rect 796 1036 804 1044
rect 844 1036 852 1044
rect 908 1036 916 1044
rect 972 1036 980 1044
rect 700 956 708 964
rect 700 936 708 944
rect 844 976 852 984
rect 892 976 900 984
rect 828 956 836 964
rect 876 956 884 964
rect 764 916 772 924
rect 796 916 804 924
rect 876 916 884 924
rect 732 896 740 904
rect 780 896 788 904
rect 892 896 900 904
rect 860 816 868 824
rect 684 776 692 784
rect 732 776 740 784
rect 300 656 308 664
rect 332 656 340 664
rect 380 656 388 664
rect 412 656 420 664
rect 284 556 292 564
rect 444 556 452 564
rect 748 556 756 564
rect 204 356 212 364
rect 316 536 324 544
rect 476 536 484 544
rect 524 536 532 544
rect 748 536 756 544
rect 572 516 580 524
rect 684 436 692 444
rect 526 406 534 414
rect 540 406 548 414
rect 554 406 562 414
rect 892 556 900 564
rect 988 916 996 924
rect 1084 896 1092 904
rect 956 816 964 824
rect 1084 816 1092 824
rect 1660 1496 1668 1504
rect 1724 1496 1732 1504
rect 1804 1502 1812 1504
rect 1804 1496 1812 1502
rect 1740 1416 1748 1424
rect 1532 1336 1540 1344
rect 1596 1336 1604 1344
rect 1660 1336 1668 1344
rect 1724 1336 1732 1344
rect 1516 1316 1524 1324
rect 1564 1316 1572 1324
rect 1596 1296 1604 1304
rect 1468 1176 1476 1184
rect 1292 1136 1300 1144
rect 1292 1116 1300 1124
rect 1548 1116 1556 1124
rect 1260 1096 1268 1104
rect 1564 1096 1572 1104
rect 1468 1076 1476 1084
rect 1260 1056 1268 1064
rect 1436 1056 1444 1064
rect 1228 1036 1236 1044
rect 1212 1016 1220 1024
rect 1148 956 1156 964
rect 1452 1036 1460 1044
rect 1420 1016 1428 1024
rect 1358 1006 1366 1014
rect 1372 1006 1380 1014
rect 1386 1006 1394 1014
rect 1372 976 1380 984
rect 1148 936 1156 944
rect 908 536 916 544
rect 732 516 740 524
rect 812 516 820 524
rect 812 436 820 444
rect 316 356 324 364
rect 428 356 436 364
rect 700 356 708 364
rect 684 336 692 344
rect 716 336 724 344
rect 252 316 260 324
rect 348 316 356 324
rect 412 316 420 324
rect 444 316 452 324
rect 588 316 596 324
rect 652 316 660 324
rect 716 316 724 324
rect 732 316 740 324
rect 252 296 260 304
rect 236 276 244 284
rect 268 276 276 284
rect 12 236 20 244
rect 44 236 52 244
rect 60 176 68 184
rect 252 256 260 264
rect 300 256 308 264
rect 204 196 212 204
rect 252 196 260 204
rect 172 136 180 144
rect 188 118 196 124
rect 188 116 196 118
rect 252 116 260 124
rect 300 176 308 184
rect 300 156 308 164
rect 412 276 420 284
rect 380 256 388 264
rect 364 236 372 244
rect 284 116 292 124
rect 316 116 324 124
rect 12 96 20 104
rect 428 176 436 184
rect 460 296 468 304
rect 524 296 532 304
rect 476 276 484 284
rect 588 276 596 284
rect 476 176 484 184
rect 796 296 804 304
rect 860 516 868 524
rect 988 696 996 704
rect 1052 696 1060 704
rect 956 656 964 664
rect 1020 676 1028 684
rect 1116 676 1124 684
rect 1004 656 1012 664
rect 972 636 980 644
rect 1052 636 1060 644
rect 1100 556 1108 564
rect 940 496 948 504
rect 844 476 852 484
rect 828 296 836 304
rect 1052 476 1060 484
rect 988 316 996 324
rect 1020 316 1028 324
rect 1164 536 1172 544
rect 1164 516 1172 524
rect 1212 936 1220 944
rect 1292 936 1300 944
rect 1340 936 1348 944
rect 1436 996 1444 1004
rect 1452 956 1460 964
rect 1436 936 1444 944
rect 1452 936 1460 944
rect 1196 916 1204 924
rect 1260 916 1268 924
rect 1308 916 1316 924
rect 1372 916 1380 924
rect 1484 956 1492 964
rect 1532 956 1540 964
rect 1676 1296 1684 1304
rect 1676 1116 1684 1124
rect 1708 1116 1716 1124
rect 1644 1096 1652 1104
rect 1628 1076 1636 1084
rect 1644 1076 1652 1084
rect 1772 1276 1780 1284
rect 1772 1256 1780 1264
rect 1884 1736 1892 1744
rect 1932 1696 1940 1704
rect 1932 1416 1940 1424
rect 1852 1256 1860 1264
rect 1772 1156 1780 1164
rect 1740 1076 1748 1084
rect 1916 1096 1924 1104
rect 1724 1036 1732 1044
rect 1708 996 1716 1004
rect 1596 976 1604 984
rect 1692 976 1700 984
rect 1516 936 1524 944
rect 1580 936 1588 944
rect 1660 936 1668 944
rect 1884 1076 1892 1084
rect 1884 1056 1892 1064
rect 1932 1056 1940 1064
rect 1804 1016 1812 1024
rect 1836 996 1844 1004
rect 1788 936 1796 944
rect 1500 916 1508 924
rect 1564 916 1572 924
rect 1644 916 1652 924
rect 1228 796 1236 804
rect 1276 796 1284 804
rect 1324 796 1332 804
rect 1532 736 1540 744
rect 1340 716 1348 724
rect 1468 716 1476 724
rect 1276 696 1284 704
rect 1388 696 1396 704
rect 1420 696 1428 704
rect 1452 696 1460 704
rect 1260 656 1268 664
rect 1292 636 1300 644
rect 1308 636 1316 644
rect 1276 576 1284 584
rect 1358 606 1366 614
rect 1372 606 1380 614
rect 1386 606 1394 614
rect 1516 656 1524 664
rect 1500 636 1508 644
rect 1452 576 1460 584
rect 1468 576 1476 584
rect 1388 556 1396 564
rect 1420 556 1428 564
rect 1436 556 1444 564
rect 1228 516 1236 524
rect 1180 456 1188 464
rect 892 296 900 304
rect 1020 296 1028 304
rect 1084 296 1092 304
rect 1132 296 1140 304
rect 1196 296 1204 304
rect 1324 496 1332 504
rect 1420 496 1428 504
rect 1484 496 1492 504
rect 844 276 852 284
rect 908 276 916 284
rect 988 276 996 284
rect 1036 276 1044 284
rect 1132 276 1140 284
rect 1164 276 1172 284
rect 1228 276 1236 284
rect 732 256 740 264
rect 396 156 404 164
rect 636 156 644 164
rect 556 136 564 144
rect 716 136 724 144
rect 780 136 788 144
rect 876 256 884 264
rect 924 256 932 264
rect 972 256 980 264
rect 1068 256 1076 264
rect 892 176 900 184
rect 924 176 932 184
rect 972 176 980 184
rect 828 136 836 144
rect 860 136 868 144
rect 380 116 388 124
rect 524 116 532 124
rect 588 118 596 124
rect 588 116 596 118
rect 636 116 644 124
rect 764 116 772 124
rect 812 116 820 124
rect 876 116 884 124
rect 1068 156 1076 164
rect 1084 136 1092 144
rect 1324 296 1332 304
rect 1388 302 1396 304
rect 1388 296 1396 302
rect 1420 296 1428 304
rect 1276 256 1284 264
rect 1292 256 1300 264
rect 1358 206 1366 214
rect 1372 206 1380 214
rect 1386 206 1394 214
rect 1164 176 1172 184
rect 1388 176 1396 184
rect 1228 156 1236 164
rect 1420 156 1428 164
rect 1548 636 1556 644
rect 1596 616 1604 624
rect 1532 596 1540 604
rect 1580 556 1588 564
rect 1580 536 1588 544
rect 1532 516 1540 524
rect 1548 496 1556 504
rect 1580 476 1588 484
rect 1916 996 1924 1004
rect 1884 976 1892 984
rect 1788 736 1796 744
rect 1660 696 1668 704
rect 1676 616 1684 624
rect 1756 616 1764 624
rect 1692 596 1700 604
rect 1740 576 1748 584
rect 1724 556 1732 564
rect 1804 556 1812 564
rect 1660 536 1668 544
rect 1804 536 1812 544
rect 1788 516 1796 524
rect 1644 476 1652 484
rect 1596 296 1604 304
rect 1516 276 1524 284
rect 1548 276 1556 284
rect 1500 136 1508 144
rect 1100 116 1108 124
rect 1164 116 1172 124
rect 1196 116 1204 124
rect 1500 116 1508 124
rect 1596 156 1604 164
rect 1596 136 1604 144
rect 1660 302 1668 304
rect 1660 296 1668 302
rect 1804 296 1812 304
rect 1788 276 1796 284
rect 1724 236 1732 244
rect 1868 896 1876 904
rect 1932 976 1940 984
rect 1836 536 1844 544
rect 1884 536 1892 544
rect 1900 516 1908 524
rect 1932 496 1940 504
rect 1836 376 1844 384
rect 1900 376 1908 384
rect 1884 276 1892 284
rect 1868 256 1876 264
rect 1644 156 1652 164
rect 1676 156 1684 164
rect 1740 156 1748 164
rect 1820 156 1828 164
rect 1900 156 1908 164
rect 1692 136 1700 144
rect 1756 136 1764 144
rect 1788 136 1796 144
rect 1852 136 1860 144
rect 1916 136 1924 144
rect 1612 116 1620 124
rect 1676 116 1684 124
rect 1724 116 1732 124
rect 1836 116 1844 124
rect 1052 96 1060 104
rect 1260 96 1268 104
rect 526 6 534 14
rect 540 6 548 14
rect 554 6 562 14
rect 1452 16 1460 24
rect 1484 16 1492 24
rect 1500 16 1508 24
rect 1532 16 1540 24
rect 1548 16 1556 24
rect 1580 16 1588 24
<< metal3 >>
rect 1352 1814 1400 1816
rect 1352 1806 1356 1814
rect 1366 1806 1372 1814
rect 1380 1806 1386 1814
rect 1396 1806 1400 1814
rect 1352 1804 1400 1806
rect 644 1797 668 1803
rect 692 1797 716 1803
rect 1860 1757 1884 1763
rect 276 1737 412 1743
rect 948 1737 1132 1743
rect 1140 1737 1468 1743
rect 1476 1737 1628 1743
rect 1636 1737 1660 1743
rect 1828 1737 1884 1743
rect 980 1717 1004 1723
rect 1716 1717 1836 1723
rect -19 1697 12 1703
rect 916 1697 1004 1703
rect 1940 1697 1971 1703
rect 13 1683 19 1696
rect 13 1677 1020 1683
rect 1316 1677 1404 1683
rect 292 1657 396 1663
rect 468 1657 700 1663
rect 740 1657 780 1663
rect 520 1614 568 1616
rect 520 1606 524 1614
rect 534 1606 540 1614
rect 548 1606 554 1614
rect 564 1606 568 1614
rect 520 1604 568 1606
rect 164 1597 236 1603
rect 244 1597 348 1603
rect 1268 1597 1292 1603
rect 596 1517 652 1523
rect 660 1517 684 1523
rect 692 1517 748 1523
rect 1236 1517 1500 1523
rect 1508 1517 1644 1523
rect 132 1497 268 1503
rect 340 1497 524 1503
rect 740 1497 828 1503
rect 836 1497 940 1503
rect 1188 1497 1260 1503
rect 1268 1497 1372 1503
rect 1396 1497 1420 1503
rect 1428 1497 1452 1503
rect 1556 1497 1660 1503
rect 1732 1497 1804 1503
rect 692 1477 716 1483
rect 820 1477 860 1483
rect 1076 1477 1164 1483
rect 1172 1477 1292 1483
rect 1300 1477 1404 1483
rect 1444 1477 1548 1483
rect 324 1457 444 1463
rect 452 1457 492 1463
rect 980 1457 1020 1463
rect 1332 1457 1436 1463
rect 1444 1457 1564 1463
rect 100 1437 204 1443
rect 212 1437 300 1443
rect 308 1437 460 1443
rect 548 1437 652 1443
rect 1380 1437 1436 1443
rect 1748 1417 1932 1423
rect 1352 1414 1400 1416
rect 1352 1406 1356 1414
rect 1366 1406 1372 1414
rect 1380 1406 1386 1414
rect 1396 1406 1400 1414
rect 1352 1404 1400 1406
rect 628 1377 844 1383
rect 1428 1377 1468 1383
rect 164 1357 204 1363
rect 260 1357 348 1363
rect 484 1357 508 1363
rect 516 1357 636 1363
rect 1204 1357 1228 1363
rect 1460 1357 1500 1363
rect 1572 1357 1612 1363
rect -19 1337 60 1343
rect 244 1337 268 1343
rect 292 1337 444 1343
rect 1012 1337 1100 1343
rect 1380 1337 1532 1343
rect 1540 1337 1596 1343
rect 1668 1337 1724 1343
rect 20 1317 44 1323
rect 52 1317 108 1323
rect 116 1317 156 1323
rect 164 1317 588 1323
rect 644 1317 732 1323
rect 804 1317 956 1323
rect 1156 1317 1228 1323
rect 1316 1317 1356 1323
rect 1364 1317 1516 1323
rect 1524 1317 1564 1323
rect -19 1297 12 1303
rect 132 1297 188 1303
rect 196 1297 364 1303
rect 692 1297 844 1303
rect 1044 1297 1276 1303
rect 1284 1297 1324 1303
rect 1604 1297 1676 1303
rect 372 1277 572 1283
rect 612 1277 636 1283
rect 644 1277 716 1283
rect 724 1277 780 1283
rect 788 1277 876 1283
rect 1268 1277 1308 1283
rect 1396 1277 1772 1283
rect 468 1257 652 1263
rect 1780 1257 1852 1263
rect 388 1237 460 1243
rect 468 1237 796 1243
rect 980 1237 988 1243
rect 520 1214 568 1216
rect 520 1206 524 1214
rect 534 1206 540 1214
rect 548 1206 554 1214
rect 564 1206 568 1214
rect 520 1204 568 1206
rect 420 1177 1196 1183
rect 1236 1177 1468 1183
rect 436 1157 620 1163
rect 628 1157 940 1163
rect 948 1157 1196 1163
rect 1204 1157 1772 1163
rect 388 1137 476 1143
rect 484 1137 588 1143
rect 596 1137 1164 1143
rect 1204 1137 1292 1143
rect 196 1117 252 1123
rect 484 1117 508 1123
rect 516 1117 636 1123
rect 708 1117 732 1123
rect 932 1117 1116 1123
rect 1268 1117 1292 1123
rect 1556 1117 1676 1123
rect 1684 1117 1708 1123
rect -19 1097 12 1103
rect 52 1097 60 1103
rect 68 1097 284 1103
rect 612 1097 652 1103
rect 740 1097 828 1103
rect 836 1097 876 1103
rect 884 1097 940 1103
rect 1108 1097 1260 1103
rect 1572 1097 1644 1103
rect 1924 1097 1971 1103
rect 228 1077 300 1083
rect 308 1077 444 1083
rect 452 1077 492 1083
rect 900 1077 956 1083
rect 1124 1077 1468 1083
rect 1476 1077 1628 1083
rect 1652 1077 1740 1083
rect 1748 1077 1884 1083
rect 292 1057 316 1063
rect 356 1057 396 1063
rect 868 1057 908 1063
rect 1268 1057 1436 1063
rect 1892 1057 1932 1063
rect 756 1037 796 1043
rect 804 1037 844 1043
rect 916 1037 972 1043
rect 1236 1037 1260 1043
rect 1460 1037 1724 1043
rect 644 1017 1212 1023
rect 1428 1017 1804 1023
rect 1352 1014 1400 1016
rect 1352 1006 1356 1014
rect 1366 1006 1372 1014
rect 1380 1006 1386 1014
rect 1396 1006 1400 1014
rect 1352 1004 1400 1006
rect 292 997 652 1003
rect 1444 997 1708 1003
rect 1716 997 1836 1003
rect 1844 997 1916 1003
rect 420 977 460 983
rect 692 977 844 983
rect 852 977 892 983
rect 1380 977 1596 983
rect 1604 977 1692 983
rect 1700 977 1884 983
rect 1940 977 1971 983
rect 132 957 252 963
rect 644 957 700 963
rect 836 957 876 963
rect 1156 957 1452 963
rect 1492 957 1532 963
rect 196 937 316 943
rect 596 937 700 943
rect 1156 937 1212 943
rect 1300 937 1340 943
rect 1348 937 1436 943
rect 1460 937 1516 943
rect 1524 937 1580 943
rect 1588 937 1660 943
rect 1796 937 1971 943
rect 100 917 364 923
rect 372 917 412 923
rect 452 917 604 923
rect 772 917 796 923
rect 884 917 988 923
rect 1204 917 1260 923
rect 1316 917 1372 923
rect 1508 917 1564 923
rect 1572 917 1644 923
rect -19 897 12 903
rect 548 897 732 903
rect 740 897 780 903
rect 788 897 892 903
rect 900 897 1084 903
rect 1876 897 1971 903
rect 308 837 364 843
rect 276 817 300 823
rect 868 817 956 823
rect 964 817 1084 823
rect 520 814 568 816
rect 520 806 524 814
rect 534 806 540 814
rect 548 806 554 814
rect 564 806 568 814
rect 520 804 568 806
rect 1236 797 1276 803
rect 1284 797 1324 803
rect 692 777 732 783
rect 1540 737 1788 743
rect 116 717 140 723
rect 180 717 204 723
rect 404 717 476 723
rect 1348 717 1468 723
rect -19 697 12 703
rect 52 697 92 703
rect 100 697 236 703
rect 244 697 316 703
rect 324 697 604 703
rect 996 697 1052 703
rect 1060 697 1276 703
rect 1396 697 1420 703
rect 1460 697 1660 703
rect 308 677 380 683
rect 1028 677 1116 683
rect 228 657 268 663
rect 276 657 300 663
rect 308 657 332 663
rect 388 657 412 663
rect 964 657 1004 663
rect 1268 657 1516 663
rect 980 637 1052 643
rect 1060 637 1292 643
rect 1300 637 1308 643
rect 1508 637 1548 643
rect 1604 617 1676 623
rect 1684 617 1756 623
rect 1352 614 1400 616
rect 1352 606 1356 614
rect 1366 606 1372 614
rect 1380 606 1386 614
rect 1396 606 1400 614
rect 1352 604 1400 606
rect 1540 597 1692 603
rect 68 577 140 583
rect 148 577 268 583
rect 1284 577 1452 583
rect 1476 577 1740 583
rect 132 557 252 563
rect 260 557 284 563
rect 452 557 748 563
rect 900 557 1100 563
rect 1396 557 1420 563
rect 1444 557 1580 563
rect 1732 557 1804 563
rect 228 537 316 543
rect 324 537 476 543
rect 484 537 524 543
rect 756 537 908 543
rect 1172 537 1580 543
rect 1588 537 1660 543
rect 1812 537 1836 543
rect 1892 537 1971 543
rect 580 517 732 523
rect 820 517 860 523
rect 1172 517 1228 523
rect 1540 517 1788 523
rect 1796 517 1900 523
rect -19 497 12 503
rect 948 497 1324 503
rect 1332 497 1420 503
rect 1492 497 1548 503
rect 1940 497 1971 503
rect 852 477 1052 483
rect 1060 477 1580 483
rect 1588 477 1644 483
rect 1188 457 1228 463
rect 692 437 812 443
rect 520 414 568 416
rect 520 406 524 414
rect 534 406 540 414
rect 548 406 554 414
rect 564 406 568 414
rect 520 404 568 406
rect 1844 377 1900 383
rect 212 357 316 363
rect 324 357 428 363
rect 436 357 700 363
rect 692 337 716 343
rect 260 317 348 323
rect 356 317 412 323
rect 452 317 588 323
rect 596 317 652 323
rect 660 317 716 323
rect 740 317 988 323
rect 1028 317 1036 323
rect 148 297 252 303
rect 468 297 524 303
rect 804 297 828 303
rect 836 297 892 303
rect 1028 297 1084 303
rect 1140 297 1196 303
rect 1332 297 1388 303
rect 1428 297 1596 303
rect 1668 297 1804 303
rect 244 277 268 283
rect 420 277 476 283
rect 596 277 844 283
rect 852 277 908 283
rect 996 277 1036 283
rect 1044 277 1132 283
rect 1172 277 1228 283
rect 1524 277 1548 283
rect 1796 277 1884 283
rect 260 257 300 263
rect 388 257 732 263
rect 884 257 924 263
rect 980 257 1068 263
rect 1204 257 1276 263
rect 1300 257 1868 263
rect 20 237 44 243
rect 52 237 364 243
rect 1277 243 1283 256
rect 1277 237 1724 243
rect 1352 214 1400 216
rect 1352 206 1356 214
rect 1366 206 1372 214
rect 1380 206 1386 214
rect 1396 206 1400 214
rect 1352 204 1400 206
rect 212 197 252 203
rect 68 177 300 183
rect 436 177 476 183
rect 900 177 924 183
rect 932 177 972 183
rect 1172 177 1388 183
rect 308 157 396 163
rect 404 157 636 163
rect 1044 157 1068 163
rect 1076 157 1228 163
rect 1236 157 1420 163
rect 1604 157 1644 163
rect 1684 157 1740 163
rect 1828 157 1900 163
rect 180 137 556 143
rect 724 137 780 143
rect 836 137 844 143
rect 868 137 1084 143
rect 1508 137 1596 143
rect 1700 137 1756 143
rect 1796 137 1852 143
rect 1860 137 1916 143
rect 196 117 252 123
rect 292 117 316 123
rect 324 117 380 123
rect 532 117 588 123
rect 644 117 764 123
rect 820 117 876 123
rect 1108 117 1164 123
rect 1204 117 1228 123
rect 1236 117 1500 123
rect 1620 117 1676 123
rect 1732 117 1836 123
rect -19 97 12 103
rect 1060 97 1260 103
rect 1460 17 1484 23
rect 1508 17 1532 23
rect 1556 17 1580 23
rect 520 14 568 16
rect 520 6 524 14
rect 534 6 540 14
rect 548 6 554 14
rect 564 6 568 14
rect 520 4 568 6
<< m4contact >>
rect 1356 1806 1358 1814
rect 1358 1806 1364 1814
rect 1372 1806 1380 1814
rect 1388 1806 1394 1814
rect 1394 1806 1396 1814
rect 972 1716 980 1724
rect 524 1606 526 1614
rect 526 1606 532 1614
rect 540 1606 548 1614
rect 556 1606 562 1614
rect 562 1606 564 1614
rect 1420 1496 1428 1504
rect 1356 1406 1358 1414
rect 1358 1406 1364 1414
rect 1372 1406 1380 1414
rect 1388 1406 1394 1414
rect 1394 1406 1396 1414
rect 1420 1376 1428 1384
rect 972 1236 980 1244
rect 524 1206 526 1214
rect 526 1206 532 1214
rect 540 1206 548 1214
rect 556 1206 562 1214
rect 562 1206 564 1214
rect 1196 1156 1204 1164
rect 1260 1116 1268 1124
rect 1260 1036 1268 1044
rect 1356 1006 1358 1014
rect 1358 1006 1364 1014
rect 1372 1006 1380 1014
rect 1388 1006 1394 1014
rect 1394 1006 1396 1014
rect 844 976 852 984
rect 524 806 526 814
rect 526 806 532 814
rect 540 806 548 814
rect 556 806 562 814
rect 562 806 564 814
rect 204 716 212 724
rect 1356 606 1358 614
rect 1358 606 1364 614
rect 1372 606 1380 614
rect 1388 606 1394 614
rect 1394 606 1396 614
rect 1228 456 1236 464
rect 524 406 526 414
rect 526 406 532 414
rect 540 406 548 414
rect 556 406 562 414
rect 562 406 564 414
rect 204 356 212 364
rect 1036 316 1044 324
rect 1196 256 1204 264
rect 1356 206 1358 214
rect 1358 206 1364 214
rect 1372 206 1380 214
rect 1388 206 1394 214
rect 1394 206 1396 214
rect 1036 156 1044 164
rect 844 136 852 144
rect 1228 116 1236 124
rect 524 6 526 14
rect 526 6 532 14
rect 540 6 548 14
rect 556 6 562 14
rect 562 6 564 14
<< metal4 >>
rect 520 1614 568 1840
rect 1352 1814 1400 1840
rect 1352 1806 1356 1814
rect 1364 1806 1372 1814
rect 1380 1806 1388 1814
rect 1396 1806 1400 1814
rect 520 1606 524 1614
rect 532 1606 540 1614
rect 548 1606 556 1614
rect 564 1606 568 1614
rect 520 1214 568 1606
rect 970 1724 982 1726
rect 970 1716 972 1724
rect 980 1716 982 1724
rect 970 1244 982 1716
rect 970 1236 972 1244
rect 980 1236 982 1244
rect 970 1234 982 1236
rect 1352 1414 1400 1806
rect 1352 1406 1356 1414
rect 1364 1406 1372 1414
rect 1380 1406 1388 1414
rect 1396 1406 1400 1414
rect 520 1206 524 1214
rect 532 1206 540 1214
rect 548 1206 556 1214
rect 564 1206 568 1214
rect 520 814 568 1206
rect 1194 1164 1206 1166
rect 1194 1156 1196 1164
rect 1204 1156 1206 1164
rect 520 806 524 814
rect 532 806 540 814
rect 548 806 556 814
rect 564 806 568 814
rect 202 724 214 726
rect 202 716 204 724
rect 212 716 214 724
rect 202 364 214 716
rect 202 356 204 364
rect 212 356 214 364
rect 202 354 214 356
rect 520 414 568 806
rect 520 406 524 414
rect 532 406 540 414
rect 548 406 556 414
rect 564 406 568 414
rect 520 14 568 406
rect 842 984 854 986
rect 842 976 844 984
rect 852 976 854 984
rect 842 144 854 976
rect 1034 324 1046 326
rect 1034 316 1036 324
rect 1044 316 1046 324
rect 1034 164 1046 316
rect 1194 264 1206 1156
rect 1258 1124 1270 1126
rect 1258 1116 1260 1124
rect 1268 1116 1270 1124
rect 1258 1044 1270 1116
rect 1258 1036 1260 1044
rect 1268 1036 1270 1044
rect 1258 1034 1270 1036
rect 1352 1014 1400 1406
rect 1418 1504 1430 1506
rect 1418 1496 1420 1504
rect 1428 1496 1430 1504
rect 1418 1384 1430 1496
rect 1418 1376 1420 1384
rect 1428 1376 1430 1384
rect 1418 1374 1430 1376
rect 1352 1006 1356 1014
rect 1364 1006 1372 1014
rect 1380 1006 1388 1014
rect 1396 1006 1400 1014
rect 1352 614 1400 1006
rect 1352 606 1356 614
rect 1364 606 1372 614
rect 1380 606 1388 614
rect 1396 606 1400 614
rect 1194 256 1196 264
rect 1204 256 1206 264
rect 1194 254 1206 256
rect 1226 464 1238 466
rect 1226 456 1228 464
rect 1236 456 1238 464
rect 1034 156 1036 164
rect 1044 156 1046 164
rect 1034 154 1046 156
rect 842 136 844 144
rect 852 136 854 144
rect 842 134 854 136
rect 1226 124 1238 456
rect 1226 116 1228 124
rect 1236 116 1238 124
rect 1226 114 1238 116
rect 1352 214 1400 606
rect 1352 206 1356 214
rect 1364 206 1372 214
rect 1380 206 1388 214
rect 1396 206 1400 214
rect 520 6 524 14
rect 532 6 540 14
rect 548 6 556 14
rect 564 6 568 14
rect 520 -40 568 6
rect 1352 -40 1400 206
use BUFX2  BUFX2_23
timestamp 1651681474
transform -1 0 56 0 -1 210
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_19
timestamp 1651681474
transform -1 0 248 0 -1 210
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_18
timestamp 1651681474
transform -1 0 200 0 1 210
box -4 -6 196 206
use OAI21X1  OAI21X1_14
timestamp 1651681474
transform -1 0 264 0 1 210
box -4 -6 68 206
use AOI21X1  AOI21X1_14
timestamp 1651681474
transform -1 0 312 0 -1 210
box -4 -6 68 206
use AND2X2  AND2X2_4
timestamp 1651681474
transform -1 0 376 0 -1 210
box -4 -6 68 206
use AOI21X1  AOI21X1_15
timestamp 1651681474
transform 1 0 376 0 -1 210
box -4 -6 68 206
use NOR2X1  NOR2X1_20
timestamp 1651681474
transform 1 0 264 0 1 210
box -4 -6 52 206
use OAI21X1  OAI21X1_13
timestamp 1651681474
transform -1 0 376 0 1 210
box -4 -6 68 206
use NAND2X1  NAND2X1_6
timestamp 1651681474
transform 1 0 376 0 1 210
box -4 -6 52 206
use NOR2X1  NOR2X1_3
timestamp 1651681474
transform 1 0 488 0 1 210
box -4 -6 52 206
use OAI21X1  OAI21X1_15
timestamp 1651681474
transform -1 0 488 0 1 210
box -4 -6 68 206
use FILL  FILL_0_0_1
timestamp 1651681474
transform 1 0 504 0 -1 210
box -4 -6 20 206
use FILL  FILL_0_0_0
timestamp 1651681474
transform 1 0 488 0 -1 210
box -4 -6 20 206
use NOR2X1  NOR2X1_21
timestamp 1651681474
transform -1 0 488 0 -1 210
box -4 -6 52 206
use NAND2X1  NAND2X1_7
timestamp 1651681474
transform -1 0 632 0 1 210
box -4 -6 52 206
use FILL  FILL_1_0_2
timestamp 1651681474
transform -1 0 584 0 1 210
box -4 -6 20 206
use FILL  FILL_1_0_1
timestamp 1651681474
transform -1 0 568 0 1 210
box -4 -6 20 206
use FILL  FILL_1_0_0
timestamp 1651681474
transform -1 0 552 0 1 210
box -4 -6 20 206
use FILL  FILL_0_0_2
timestamp 1651681474
transform 1 0 520 0 -1 210
box -4 -6 20 206
use DFFPOSX1  DFFPOSX1_20
timestamp 1651681474
transform 1 0 536 0 -1 210
box -4 -6 196 206
use BUFX2  BUFX2_24
timestamp 1651681474
transform -1 0 776 0 -1 210
box -4 -6 52 206
use BUFX2  BUFX2_25
timestamp 1651681474
transform 1 0 776 0 -1 210
box -4 -6 52 206
use AND2X2  AND2X2_5
timestamp 1651681474
transform 1 0 632 0 1 210
box -4 -6 68 206
use NAND3X1  NAND3X1_1
timestamp 1651681474
transform -1 0 760 0 1 210
box -4 -6 68 206
use AND2X2  AND2X2_3
timestamp 1651681474
transform -1 0 824 0 1 210
box -4 -6 68 206
use BUFX2  BUFX2_20
timestamp 1651681474
transform 1 0 824 0 -1 210
box -4 -6 52 206
use BUFX2  BUFX2_27
timestamp 1651681474
transform 1 0 872 0 -1 210
box -4 -6 52 206
use BUFX2  BUFX2_26
timestamp 1651681474
transform 1 0 920 0 -1 210
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_21
timestamp 1651681474
transform -1 0 1160 0 -1 210
box -4 -6 196 206
use AOI21X1  AOI21X1_16
timestamp 1651681474
transform 1 0 824 0 1 210
box -4 -6 68 206
use OAI21X1  OAI21X1_16
timestamp 1651681474
transform 1 0 888 0 1 210
box -4 -6 68 206
use OAI21X1  OAI21X1_17
timestamp 1651681474
transform -1 0 1016 0 1 210
box -4 -6 68 206
use NAND2X1  NAND2X1_2
timestamp 1651681474
transform -1 0 1208 0 -1 210
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_23
timestamp 1651681474
transform 1 0 1208 0 -1 210
box -4 -6 196 206
use AOI21X1  AOI21X1_18
timestamp 1651681474
transform 1 0 1016 0 1 210
box -4 -6 68 206
use INVX1  INVX1_14
timestamp 1651681474
transform -1 0 1112 0 1 210
box -4 -6 36 206
use OAI21X1  OAI21X1_18
timestamp 1651681474
transform 1 0 1112 0 1 210
box -4 -6 68 206
use OAI21X1  OAI21X1_19
timestamp 1651681474
transform 1 0 1176 0 1 210
box -4 -6 68 206
use FILL  FILL_0_1_0
timestamp 1651681474
transform 1 0 1400 0 -1 210
box -4 -6 20 206
use NOR2X1  NOR2X1_23
timestamp 1651681474
transform -1 0 1288 0 1 210
box -4 -6 52 206
use FILL  FILL_1_1_0
timestamp 1651681474
transform 1 0 1288 0 1 210
box -4 -6 20 206
use FILL  FILL_1_1_1
timestamp 1651681474
transform 1 0 1304 0 1 210
box -4 -6 20 206
use FILL  FILL_1_1_2
timestamp 1651681474
transform 1 0 1320 0 1 210
box -4 -6 20 206
use DFFPOSX1  DFFPOSX1_24
timestamp 1651681474
transform 1 0 1336 0 1 210
box -4 -6 196 206
use FILL  FILL_0_1_1
timestamp 1651681474
transform 1 0 1416 0 -1 210
box -4 -6 20 206
use FILL  FILL_0_1_2
timestamp 1651681474
transform 1 0 1432 0 -1 210
box -4 -6 20 206
use BUFX2  BUFX2_28
timestamp 1651681474
transform 1 0 1448 0 -1 210
box -4 -6 52 206
use BUFX2  BUFX2_29
timestamp 1651681474
transform 1 0 1496 0 -1 210
box -4 -6 52 206
use BUFX2  BUFX2_30
timestamp 1651681474
transform 1 0 1544 0 -1 210
box -4 -6 52 206
use BUFX2  BUFX2_31
timestamp 1651681474
transform 1 0 1592 0 -1 210
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_27
timestamp 1651681474
transform -1 0 1720 0 1 210
box -4 -6 196 206
use INVX1  INVX1_18
timestamp 1651681474
transform 1 0 1640 0 -1 210
box -4 -6 36 206
use AOI21X1  AOI21X1_20
timestamp 1651681474
transform 1 0 1672 0 -1 210
box -4 -6 68 206
use OR2X2  OR2X2_4
timestamp 1651681474
transform 1 0 1736 0 -1 210
box -4 -6 68 206
use AND2X2  AND2X2_14
timestamp 1651681474
transform -1 0 1864 0 -1 210
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_28
timestamp 1651681474
transform 1 0 1720 0 1 210
box -4 -6 196 206
use AOI21X1  AOI21X1_21
timestamp 1651681474
transform -1 0 1928 0 -1 210
box -4 -6 68 206
use FILL  FILL_1_1
timestamp 1651681474
transform -1 0 1944 0 -1 210
box -4 -6 20 206
use FILL  FILL_2_1
timestamp 1651681474
transform 1 0 1912 0 1 210
box -4 -6 20 206
use FILL  FILL_2_2
timestamp 1651681474
transform 1 0 1928 0 1 210
box -4 -6 20 206
use BUFX2  BUFX2_7
timestamp 1651681474
transform -1 0 56 0 -1 610
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_2
timestamp 1651681474
transform -1 0 248 0 -1 610
box -4 -6 196 206
use AND2X2  AND2X2_7
timestamp 1651681474
transform 1 0 248 0 -1 610
box -4 -6 68 206
use CLKBUF1  CLKBUF1_3
timestamp 1651681474
transform -1 0 456 0 -1 610
box -4 -6 148 206
use FILL  FILL_2_0_0
timestamp 1651681474
transform 1 0 456 0 -1 610
box -4 -6 20 206
use FILL  FILL_2_0_1
timestamp 1651681474
transform 1 0 472 0 -1 610
box -4 -6 20 206
use FILL  FILL_2_0_2
timestamp 1651681474
transform 1 0 488 0 -1 610
box -4 -6 20 206
use DFFPOSX1  DFFPOSX1_22
timestamp 1651681474
transform 1 0 504 0 -1 610
box -4 -6 196 206
use NAND2X1  NAND2X1_21
timestamp 1651681474
transform 1 0 696 0 -1 610
box -4 -6 52 206
use NOR2X1  NOR2X1_22
timestamp 1651681474
transform 1 0 744 0 -1 610
box -4 -6 52 206
use AOI21X1  AOI21X1_17
timestamp 1651681474
transform -1 0 856 0 -1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_5
timestamp 1651681474
transform 1 0 856 0 -1 610
box -4 -6 52 206
use CLKBUF1  CLKBUF1_2
timestamp 1651681474
transform 1 0 904 0 -1 610
box -4 -6 148 206
use NAND2X1  NAND2X1_22
timestamp 1651681474
transform -1 0 1096 0 -1 610
box -4 -6 52 206
use NOR2X1  NOR2X1_2
timestamp 1651681474
transform 1 0 1096 0 -1 610
box -4 -6 52 206
use NOR3X1  NOR3X1_1
timestamp 1651681474
transform -1 0 1272 0 -1 610
box -4 -6 132 206
use OAI21X1  OAI21X1_22
timestamp 1651681474
transform 1 0 1272 0 -1 610
box -4 -6 68 206
use FILL  FILL_2_1_0
timestamp 1651681474
transform -1 0 1352 0 -1 610
box -4 -6 20 206
use FILL  FILL_2_1_1
timestamp 1651681474
transform -1 0 1368 0 -1 610
box -4 -6 20 206
use FILL  FILL_2_1_2
timestamp 1651681474
transform -1 0 1384 0 -1 610
box -4 -6 20 206
use AND2X2  AND2X2_12
timestamp 1651681474
transform -1 0 1448 0 -1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_1
timestamp 1651681474
transform -1 0 1496 0 -1 610
box -4 -6 52 206
use AND2X2  AND2X2_1
timestamp 1651681474
transform 1 0 1496 0 -1 610
box -4 -6 68 206
use NAND3X1  NAND3X1_8
timestamp 1651681474
transform 1 0 1560 0 -1 610
box -4 -6 68 206
use NAND3X1  NAND3X1_3
timestamp 1651681474
transform -1 0 1688 0 -1 610
box -4 -6 68 206
use NOR2X1  NOR2X1_1
timestamp 1651681474
transform 1 0 1688 0 -1 610
box -4 -6 52 206
use AND2X2  AND2X2_2
timestamp 1651681474
transform -1 0 1800 0 -1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_4
timestamp 1651681474
transform -1 0 1848 0 -1 610
box -4 -6 52 206
use BUFX2  BUFX2_33
timestamp 1651681474
transform 1 0 1848 0 -1 610
box -4 -6 52 206
use BUFX2  BUFX2_32
timestamp 1651681474
transform 1 0 1896 0 -1 610
box -4 -6 52 206
use BUFX2  BUFX2_8
timestamp 1651681474
transform -1 0 56 0 1 610
box -4 -6 52 206
use NAND3X1  NAND3X1_5
timestamp 1651681474
transform -1 0 120 0 1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_3
timestamp 1651681474
transform 1 0 120 0 1 610
box -4 -6 68 206
use NOR2X1  NOR2X1_5
timestamp 1651681474
transform -1 0 232 0 1 610
box -4 -6 52 206
use NAND2X1  NAND2X1_9
timestamp 1651681474
transform 1 0 232 0 1 610
box -4 -6 52 206
use INVX1  INVX1_4
timestamp 1651681474
transform 1 0 280 0 1 610
box -4 -6 36 206
use OAI21X1  OAI21X1_4
timestamp 1651681474
transform 1 0 312 0 1 610
box -4 -6 68 206
use NOR2X1  NOR2X1_6
timestamp 1651681474
transform -1 0 424 0 1 610
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_3
timestamp 1651681474
transform 1 0 424 0 1 610
box -4 -6 196 206
use FILL  FILL_3_0_0
timestamp 1651681474
transform 1 0 616 0 1 610
box -4 -6 20 206
use FILL  FILL_3_0_1
timestamp 1651681474
transform 1 0 632 0 1 610
box -4 -6 20 206
use FILL  FILL_3_0_2
timestamp 1651681474
transform 1 0 648 0 1 610
box -4 -6 20 206
use INVX1  INVX1_2
timestamp 1651681474
transform 1 0 664 0 1 610
box -4 -6 36 206
use BUFX2  BUFX2_3
timestamp 1651681474
transform -1 0 744 0 1 610
box -4 -6 52 206
use CLKBUF1  CLKBUF1_1
timestamp 1651681474
transform 1 0 744 0 1 610
box -4 -6 148 206
use BUFX2  BUFX2_4
timestamp 1651681474
transform 1 0 888 0 1 610
box -4 -6 52 206
use OAI21X1  OAI21X1_20
timestamp 1651681474
transform -1 0 1000 0 1 610
box -4 -6 68 206
use AOI21X1  AOI21X1_19
timestamp 1651681474
transform -1 0 1064 0 1 610
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_25
timestamp 1651681474
transform 1 0 1064 0 1 610
box -4 -6 196 206
use INVX1  INVX1_16
timestamp 1651681474
transform 1 0 1256 0 1 610
box -4 -6 36 206
use OAI21X1  OAI21X1_21
timestamp 1651681474
transform 1 0 1288 0 1 610
box -4 -6 68 206
use FILL  FILL_3_1_0
timestamp 1651681474
transform 1 0 1352 0 1 610
box -4 -6 20 206
use FILL  FILL_3_1_1
timestamp 1651681474
transform 1 0 1368 0 1 610
box -4 -6 20 206
use FILL  FILL_3_1_2
timestamp 1651681474
transform 1 0 1384 0 1 610
box -4 -6 20 206
use AND2X2  AND2X2_13
timestamp 1651681474
transform 1 0 1400 0 1 610
box -4 -6 68 206
use INVX1  INVX1_17
timestamp 1651681474
transform -1 0 1496 0 1 610
box -4 -6 36 206
use NAND2X1  NAND2X1_3
timestamp 1651681474
transform 1 0 1496 0 1 610
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_26
timestamp 1651681474
transform -1 0 1736 0 1 610
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_29
timestamp 1651681474
transform 1 0 1736 0 1 610
box -4 -6 196 206
use FILL  FILL_4_1
timestamp 1651681474
transform 1 0 1928 0 1 610
box -4 -6 20 206
use BUFX2  BUFX2_9
timestamp 1651681474
transform -1 0 56 0 -1 1010
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_4
timestamp 1651681474
transform -1 0 248 0 -1 1010
box -4 -6 196 206
use OAI21X1  OAI21X1_5
timestamp 1651681474
transform 1 0 248 0 -1 1010
box -4 -6 68 206
use NOR2X1  NOR2X1_8
timestamp 1651681474
transform -1 0 360 0 -1 1010
box -4 -6 52 206
use NOR2X1  NOR2X1_7
timestamp 1651681474
transform -1 0 408 0 -1 1010
box -4 -6 52 206
use INVX1  INVX1_7
timestamp 1651681474
transform 1 0 408 0 -1 1010
box -4 -6 36 206
use NAND2X1  NAND2X1_12
timestamp 1651681474
transform 1 0 440 0 -1 1010
box -4 -6 52 206
use BUFX2  BUFX2_2
timestamp 1651681474
transform -1 0 536 0 -1 1010
box -4 -6 52 206
use FILL  FILL_4_0_0
timestamp 1651681474
transform 1 0 536 0 -1 1010
box -4 -6 20 206
use FILL  FILL_4_0_1
timestamp 1651681474
transform 1 0 552 0 -1 1010
box -4 -6 20 206
use FILL  FILL_4_0_2
timestamp 1651681474
transform 1 0 568 0 -1 1010
box -4 -6 20 206
use AND2X2  AND2X2_10
timestamp 1651681474
transform 1 0 584 0 -1 1010
box -4 -6 68 206
use NAND2X1  NAND2X1_18
timestamp 1651681474
transform 1 0 648 0 -1 1010
box -4 -6 52 206
use NOR2X1  NOR2X1_18
timestamp 1651681474
transform -1 0 744 0 -1 1010
box -4 -6 52 206
use BUFX2  BUFX2_5
timestamp 1651681474
transform -1 0 792 0 -1 1010
box -4 -6 52 206
use NOR2X1  NOR2X1_17
timestamp 1651681474
transform -1 0 840 0 -1 1010
box -4 -6 52 206
use NOR2X1  NOR2X1_19
timestamp 1651681474
transform -1 0 888 0 -1 1010
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_15
timestamp 1651681474
transform -1 0 1080 0 -1 1010
box -4 -6 196 206
use BUFX2  BUFX2_1
timestamp 1651681474
transform 1 0 1080 0 -1 1010
box -4 -6 52 206
use INVX1  INVX1_1
timestamp 1651681474
transform -1 0 1160 0 -1 1010
box -4 -6 36 206
use INVX1  INVX1_15
timestamp 1651681474
transform -1 0 1192 0 -1 1010
box -4 -6 36 206
use AOI21X1  AOI21X1_1
timestamp 1651681474
transform 1 0 1192 0 -1 1010
box -4 -6 68 206
use NAND3X1  NAND3X1_2
timestamp 1651681474
transform -1 0 1320 0 -1 1010
box -4 -6 68 206
use AOI21X1  AOI21X1_23
timestamp 1651681474
transform 1 0 1320 0 -1 1010
box -4 -6 68 206
use FILL  FILL_4_1_0
timestamp 1651681474
transform 1 0 1384 0 -1 1010
box -4 -6 20 206
use FILL  FILL_4_1_1
timestamp 1651681474
transform 1 0 1400 0 -1 1010
box -4 -6 20 206
use FILL  FILL_4_1_2
timestamp 1651681474
transform 1 0 1416 0 -1 1010
box -4 -6 20 206
use INVX1  INVX1_20
timestamp 1651681474
transform 1 0 1432 0 -1 1010
box -4 -6 36 206
use OAI21X1  OAI21X1_23
timestamp 1651681474
transform -1 0 1528 0 -1 1010
box -4 -6 68 206
use AOI21X1  AOI21X1_22
timestamp 1651681474
transform -1 0 1592 0 -1 1010
box -4 -6 68 206
use INVX1  INVX1_21
timestamp 1651681474
transform 1 0 1592 0 -1 1010
box -4 -6 36 206
use NOR3X1  NOR3X1_2
timestamp 1651681474
transform 1 0 1624 0 -1 1010
box -4 -6 132 206
use BUFX2  BUFX2_36
timestamp 1651681474
transform 1 0 1752 0 -1 1010
box -4 -6 52 206
use INVX1  INVX1_19
timestamp 1651681474
transform -1 0 1832 0 -1 1010
box -4 -6 36 206
use BUFX2  BUFX2_34
timestamp 1651681474
transform 1 0 1832 0 -1 1010
box -4 -6 52 206
use BUFX2  BUFX2_35
timestamp 1651681474
transform 1 0 1880 0 -1 1010
box -4 -6 52 206
use FILL  FILL_5_1
timestamp 1651681474
transform -1 0 1944 0 -1 1010
box -4 -6 20 206
use BUFX2  BUFX2_6
timestamp 1651681474
transform -1 0 56 0 1 1010
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_1
timestamp 1651681474
transform -1 0 248 0 1 1010
box -4 -6 196 206
use AND2X2  AND2X2_6
timestamp 1651681474
transform -1 0 312 0 1 1010
box -4 -6 68 206
use INVX1  INVX1_5
timestamp 1651681474
transform 1 0 312 0 1 1010
box -4 -6 36 206
use NOR2X1  NOR2X1_13
timestamp 1651681474
transform 1 0 344 0 1 1010
box -4 -6 52 206
use OAI21X1  OAI21X1_9
timestamp 1651681474
transform 1 0 392 0 1 1010
box -4 -6 68 206
use NAND3X1  NAND3X1_6
timestamp 1651681474
transform -1 0 520 0 1 1010
box -4 -6 68 206
use FILL  FILL_5_0_0
timestamp 1651681474
transform -1 0 536 0 1 1010
box -4 -6 20 206
use FILL  FILL_5_0_1
timestamp 1651681474
transform -1 0 552 0 1 1010
box -4 -6 20 206
use FILL  FILL_5_0_2
timestamp 1651681474
transform -1 0 568 0 1 1010
box -4 -6 20 206
use NAND3X1  NAND3X1_7
timestamp 1651681474
transform -1 0 632 0 1 1010
box -4 -6 68 206
use AND2X2  AND2X2_11
timestamp 1651681474
transform 1 0 632 0 1 1010
box -4 -6 68 206
use NAND2X1  NAND2X1_19
timestamp 1651681474
transform 1 0 696 0 1 1010
box -4 -6 52 206
use NOR2X1  NOR2X1_16
timestamp 1651681474
transform 1 0 744 0 1 1010
box -4 -6 52 206
use NAND2X1  NAND2X1_20
timestamp 1651681474
transform 1 0 792 0 1 1010
box -4 -6 52 206
use OAI21X1  OAI21X1_12
timestamp 1651681474
transform -1 0 904 0 1 1010
box -4 -6 68 206
use AOI21X1  AOI21X1_13
timestamp 1651681474
transform -1 0 968 0 1 1010
box -4 -6 68 206
use INVX1  INVX1_13
timestamp 1651681474
transform -1 0 1000 0 1 1010
box -4 -6 36 206
use DFFPOSX1  DFFPOSX1_16
timestamp 1651681474
transform -1 0 1192 0 1 1010
box -4 -6 196 206
use NOR2X1  NOR2X1_11
timestamp 1651681474
transform -1 0 1240 0 1 1010
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_31
timestamp 1651681474
transform 1 0 1240 0 1 1010
box -4 -6 196 206
use FILL  FILL_5_1_0
timestamp 1651681474
transform -1 0 1448 0 1 1010
box -4 -6 20 206
use FILL  FILL_5_1_1
timestamp 1651681474
transform -1 0 1464 0 1 1010
box -4 -6 20 206
use FILL  FILL_5_1_2
timestamp 1651681474
transform -1 0 1480 0 1 1010
box -4 -6 20 206
use OAI21X1  OAI21X1_1
timestamp 1651681474
transform -1 0 1544 0 1 1010
box -4 -6 68 206
use OAI21X1  OAI21X1_2
timestamp 1651681474
transform 1 0 1544 0 1 1010
box -4 -6 68 206
use INVX1  INVX1_3
timestamp 1651681474
transform -1 0 1640 0 1 1010
box -4 -6 36 206
use NOR2X1  NOR2X1_4
timestamp 1651681474
transform -1 0 1688 0 1 1010
box -4 -6 52 206
use NAND3X1  NAND3X1_4
timestamp 1651681474
transform 1 0 1688 0 1 1010
box -4 -6 68 206
use NOR3X1  NOR3X1_3
timestamp 1651681474
transform 1 0 1752 0 1 1010
box -4 -6 132 206
use BUFX2  BUFX2_37
timestamp 1651681474
transform 1 0 1880 0 1 1010
box -4 -6 52 206
use FILL  FILL_6_1
timestamp 1651681474
transform 1 0 1928 0 1 1010
box -4 -6 20 206
use BUFX2  BUFX2_14
timestamp 1651681474
transform -1 0 56 0 -1 1410
box -4 -6 52 206
use BUFX2  BUFX2_17
timestamp 1651681474
transform -1 0 104 0 -1 1410
box -4 -6 52 206
use AOI21X1  AOI21X1_7
timestamp 1651681474
transform 1 0 104 0 -1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_10
timestamp 1651681474
transform 1 0 168 0 -1 1410
box -4 -6 68 206
use INVX1  INVX1_9
timestamp 1651681474
transform 1 0 232 0 -1 1410
box -4 -6 36 206
use NAND2X1  NAND2X1_15
timestamp 1651681474
transform 1 0 264 0 -1 1410
box -4 -6 52 206
use OR2X2  OR2X2_1
timestamp 1651681474
transform -1 0 376 0 -1 1410
box -4 -6 68 206
use AOI21X1  AOI21X1_9
timestamp 1651681474
transform 1 0 376 0 -1 1410
box -4 -6 68 206
use NOR2X1  NOR2X1_15
timestamp 1651681474
transform -1 0 488 0 -1 1410
box -4 -6 52 206
use INVX1  INVX1_8
timestamp 1651681474
transform -1 0 520 0 -1 1410
box -4 -6 36 206
use FILL  FILL_6_0_0
timestamp 1651681474
transform 1 0 520 0 -1 1410
box -4 -6 20 206
use FILL  FILL_6_0_1
timestamp 1651681474
transform 1 0 536 0 -1 1410
box -4 -6 20 206
use FILL  FILL_6_0_2
timestamp 1651681474
transform 1 0 552 0 -1 1410
box -4 -6 20 206
use AOI21X1  AOI21X1_8
timestamp 1651681474
transform 1 0 568 0 -1 1410
box -4 -6 68 206
use NAND2X1  NAND2X1_16
timestamp 1651681474
transform -1 0 680 0 -1 1410
box -4 -6 52 206
use OAI21X1  OAI21X1_11
timestamp 1651681474
transform -1 0 744 0 -1 1410
box -4 -6 68 206
use NOR2X1  NOR2X1_14
timestamp 1651681474
transform -1 0 792 0 -1 1410
box -4 -6 52 206
use NAND2X1  NAND2X1_14
timestamp 1651681474
transform -1 0 840 0 -1 1410
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_10
timestamp 1651681474
transform -1 0 1032 0 -1 1410
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_8
timestamp 1651681474
transform -1 0 1224 0 -1 1410
box -4 -6 196 206
use NOR2X1  NOR2X1_12
timestamp 1651681474
transform 1 0 1224 0 -1 1410
box -4 -6 52 206
use NAND2X1  NAND2X1_11
timestamp 1651681474
transform -1 0 1320 0 -1 1410
box -4 -6 52 206
use AOI21X1  AOI21X1_6
timestamp 1651681474
transform -1 0 1384 0 -1 1410
box -4 -6 68 206
use FILL  FILL_6_1_0
timestamp 1651681474
transform 1 0 1384 0 -1 1410
box -4 -6 20 206
use FILL  FILL_6_1_1
timestamp 1651681474
transform 1 0 1400 0 -1 1410
box -4 -6 20 206
use FILL  FILL_6_1_2
timestamp 1651681474
transform 1 0 1416 0 -1 1410
box -4 -6 20 206
use INVX1  INVX1_6
timestamp 1651681474
transform 1 0 1432 0 -1 1410
box -4 -6 36 206
use NOR2X1  NOR2X1_10
timestamp 1651681474
transform 1 0 1464 0 -1 1410
box -4 -6 52 206
use AOI21X1  AOI21X1_5
timestamp 1651681474
transform 1 0 1512 0 -1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_8
timestamp 1651681474
transform 1 0 1576 0 -1 1410
box -4 -6 68 206
use NAND2X1  NAND2X1_8
timestamp 1651681474
transform 1 0 1640 0 -1 1410
box -4 -6 52 206
use AOI21X1  AOI21X1_2
timestamp 1651681474
transform -1 0 1752 0 -1 1410
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_30
timestamp 1651681474
transform 1 0 1752 0 -1 1410
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_9
timestamp 1651681474
transform -1 0 200 0 1 1410
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_12
timestamp 1651681474
transform -1 0 392 0 1 1410
box -4 -6 196 206
use AND2X2  AND2X2_8
timestamp 1651681474
transform -1 0 456 0 1 1410
box -4 -6 68 206
use INVX1  INVX1_10
timestamp 1651681474
transform 1 0 456 0 1 1410
box -4 -6 36 206
use AOI21X1  AOI21X1_10
timestamp 1651681474
transform 1 0 488 0 1 1410
box -4 -6 68 206
use FILL  FILL_7_0_0
timestamp 1651681474
transform 1 0 552 0 1 1410
box -4 -6 20 206
use FILL  FILL_7_0_1
timestamp 1651681474
transform 1 0 568 0 1 1410
box -4 -6 20 206
use FILL  FILL_7_0_2
timestamp 1651681474
transform 1 0 584 0 1 1410
box -4 -6 20 206
use NAND2X1  NAND2X1_13
timestamp 1651681474
transform 1 0 600 0 1 1410
box -4 -6 52 206
use INVX1  INVX1_12
timestamp 1651681474
transform 1 0 648 0 1 1410
box -4 -6 36 206
use AOI21X1  AOI21X1_12
timestamp 1651681474
transform -1 0 744 0 1 1410
box -4 -6 68 206
use NAND2X1  NAND2X1_17
timestamp 1651681474
transform -1 0 792 0 1 1410
box -4 -6 52 206
use INVX1  INVX1_11
timestamp 1651681474
transform 1 0 792 0 1 1410
box -4 -6 36 206
use OR2X2  OR2X2_2
timestamp 1651681474
transform -1 0 888 0 1 1410
box -4 -6 68 206
use AOI21X1  AOI21X1_11
timestamp 1651681474
transform 1 0 888 0 1 1410
box -4 -6 68 206
use AND2X2  AND2X2_9
timestamp 1651681474
transform 1 0 952 0 1 1410
box -4 -6 68 206
use CLKBUF1  CLKBUF1_5
timestamp 1651681474
transform 1 0 1016 0 1 1410
box -4 -6 148 206
use AOI21X1  AOI21X1_3
timestamp 1651681474
transform 1 0 1160 0 1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_6
timestamp 1651681474
transform -1 0 1288 0 1 1410
box -4 -6 68 206
use NAND2X1  NAND2X1_10
timestamp 1651681474
transform 1 0 1288 0 1 1410
box -4 -6 52 206
use FILL  FILL_7_1_0
timestamp 1651681474
transform 1 0 1336 0 1 1410
box -4 -6 20 206
use FILL  FILL_7_1_1
timestamp 1651681474
transform 1 0 1352 0 1 1410
box -4 -6 20 206
use FILL  FILL_7_1_2
timestamp 1651681474
transform 1 0 1368 0 1 1410
box -4 -6 20 206
use AOI21X1  AOI21X1_4
timestamp 1651681474
transform 1 0 1384 0 1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_7
timestamp 1651681474
transform 1 0 1448 0 1 1410
box -4 -6 68 206
use NOR2X1  NOR2X1_9
timestamp 1651681474
transform -1 0 1560 0 1 1410
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_6
timestamp 1651681474
transform -1 0 1752 0 1 1410
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_32
timestamp 1651681474
transform 1 0 1752 0 1 1410
box -4 -6 196 206
use CLKBUF1  CLKBUF1_4
timestamp 1651681474
transform 1 0 8 0 -1 1810
box -4 -6 148 206
use DFFPOSX1  DFFPOSX1_11
timestamp 1651681474
transform -1 0 344 0 -1 1810
box -4 -6 196 206
use BUFX2  BUFX2_16
timestamp 1651681474
transform 1 0 344 0 -1 1810
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_14
timestamp 1651681474
transform 1 0 392 0 -1 1810
box -4 -6 196 206
use FILL  FILL_8_0_0
timestamp 1651681474
transform 1 0 584 0 -1 1810
box -4 -6 20 206
use FILL  FILL_8_0_1
timestamp 1651681474
transform 1 0 600 0 -1 1810
box -4 -6 20 206
use FILL  FILL_8_0_2
timestamp 1651681474
transform 1 0 616 0 -1 1810
box -4 -6 20 206
use BUFX2  BUFX2_15
timestamp 1651681474
transform 1 0 632 0 -1 1810
box -4 -6 52 206
use BUFX2  BUFX2_19
timestamp 1651681474
transform 1 0 680 0 -1 1810
box -4 -6 52 206
use BUFX2  BUFX2_18
timestamp 1651681474
transform 1 0 728 0 -1 1810
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_13
timestamp 1651681474
transform -1 0 968 0 -1 1810
box -4 -6 196 206
use BUFX2  BUFX2_21
timestamp 1651681474
transform -1 0 1016 0 -1 1810
box -4 -6 52 206
use BUFX2  BUFX2_13
timestamp 1651681474
transform -1 0 1064 0 -1 1810
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_5
timestamp 1651681474
transform -1 0 1256 0 -1 1810
box -4 -6 196 206
use BUFX2  BUFX2_10
timestamp 1651681474
transform 1 0 1256 0 -1 1810
box -4 -6 52 206
use BUFX2  BUFX2_12
timestamp 1651681474
transform 1 0 1304 0 -1 1810
box -4 -6 52 206
use FILL  FILL_8_1_0
timestamp 1651681474
transform -1 0 1368 0 -1 1810
box -4 -6 20 206
use FILL  FILL_8_1_1
timestamp 1651681474
transform -1 0 1384 0 -1 1810
box -4 -6 20 206
use FILL  FILL_8_1_2
timestamp 1651681474
transform -1 0 1400 0 -1 1810
box -4 -6 20 206
use DFFPOSX1  DFFPOSX1_7
timestamp 1651681474
transform -1 0 1592 0 -1 1810
box -4 -6 196 206
use BUFX2  BUFX2_11
timestamp 1651681474
transform 1 0 1592 0 -1 1810
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_17
timestamp 1651681474
transform 1 0 1640 0 -1 1810
box -4 -6 196 206
use OR2X2  OR2X2_3
timestamp 1651681474
transform -1 0 1896 0 -1 1810
box -4 -6 68 206
use BUFX2  BUFX2_22
timestamp 1651681474
transform 1 0 1896 0 -1 1810
box -4 -6 52 206
<< labels >>
flabel metal4 s 520 -40 568 -16 7 FreeSans 24 270 0 0 vdd
port 0 nsew
flabel metal4 s 1352 -40 1400 -16 7 FreeSans 24 270 0 0 gnd
port 1 nsew
flabel metal2 s 333 -23 339 -17 7 FreeSans 24 270 0 0 address_enable
port 2 nsew
flabel metal3 s -19 1697 -13 1703 7 FreeSans 24 0 0 0 clock
port 3 nsew
flabel metal2 s 1853 1837 1859 1843 3 FreeSans 24 90 0 0 reset
port 4 nsew
flabel metal3 s -19 1097 -13 1103 7 FreeSans 24 0 0 0 address_a[0]
port 5 nsew
flabel metal3 s -19 497 -13 503 7 FreeSans 24 0 0 0 address_a[1]
port 6 nsew
flabel metal3 s -19 697 -13 703 7 FreeSans 24 0 0 0 address_a[2]
port 7 nsew
flabel metal3 s -19 897 -13 903 7 FreeSans 24 0 0 0 address_a[3]
port 8 nsew
flabel metal2 s 1277 1837 1283 1843 3 FreeSans 24 90 0 0 address_a[4]
port 9 nsew
flabel metal2 s 1613 1837 1619 1843 3 FreeSans 24 90 0 0 address_a[5]
port 10 nsew
flabel metal2 s 1325 1837 1331 1843 3 FreeSans 24 90 0 0 address_a[6]
port 11 nsew
flabel metal2 s 1037 1837 1043 1843 3 FreeSans 24 90 0 0 address_a[7]
port 12 nsew
flabel metal3 s -19 1297 -13 1303 7 FreeSans 24 0 0 0 address_a[8]
port 13 nsew
flabel metal2 s 637 1837 643 1843 3 FreeSans 24 90 0 0 address_a[9]
port 14 nsew
flabel metal2 s 365 1837 371 1843 3 FreeSans 24 90 0 0 address_a[10]
port 15 nsew
flabel metal3 s -19 1337 -13 1343 7 FreeSans 24 0 0 0 address_a[11]
port 16 nsew
flabel metal2 s 749 1837 755 1843 3 FreeSans 24 90 0 0 address_a[12]
port 17 nsew
flabel metal2 s 685 1837 691 1843 3 FreeSans 24 90 0 0 address_a[13]
port 18 nsew
flabel metal2 s 845 -23 851 -17 7 FreeSans 24 270 0 0 address_a[14]
port 19 nsew
flabel metal2 s 989 1837 995 1843 3 FreeSans 24 90 0 0 address_a[15]
port 20 nsew
flabel metal3 s 1965 1697 1971 1703 3 FreeSans 24 0 0 0 address_b[0]
port 21 nsew
flabel metal3 s -19 97 -13 103 7 FreeSans 24 0 0 0 address_b[1]
port 22 nsew
flabel metal2 s 733 -23 739 -17 7 FreeSans 24 270 0 0 address_b[2]
port 23 nsew
flabel metal2 s 797 -23 803 -17 7 FreeSans 24 270 0 0 address_b[3]
port 24 nsew
flabel metal2 s 941 -23 947 -17 7 FreeSans 24 270 0 0 address_b[4]
port 25 nsew
flabel metal2 s 893 -23 899 -17 7 FreeSans 24 270 0 0 address_b[5]
port 26 nsew
flabel metal2 s 1453 -23 1459 -17 7 FreeSans 24 270 0 0 address_b[6]
port 27 nsew
flabel metal2 s 1501 -23 1507 -17 7 FreeSans 24 270 0 0 address_b[7]
port 28 nsew
flabel metal2 s 1549 -23 1555 -17 7 FreeSans 24 270 0 0 address_b[8]
port 29 nsew
flabel metal2 s 1613 -23 1619 -17 7 FreeSans 24 270 0 0 address_b[9]
port 30 nsew
flabel metal3 s 1965 497 1971 503 3 FreeSans 24 0 0 0 address_b[10]
port 31 nsew
flabel metal3 s 1965 537 1971 543 3 FreeSans 24 0 0 0 address_b[11]
port 32 nsew
flabel metal3 s 1965 897 1971 903 3 FreeSans 24 0 0 0 address_b[12]
port 33 nsew
flabel metal3 s 1965 977 1971 983 3 FreeSans 24 0 0 0 address_b[13]
port 34 nsew
flabel metal3 s 1965 937 1971 943 3 FreeSans 24 0 0 0 address_b[14]
port 35 nsew
flabel metal3 s 1965 1097 1971 1103 3 FreeSans 24 0 0 0 address_b[15]
port 36 nsew
<< end >>
