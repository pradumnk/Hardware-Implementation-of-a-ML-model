magic
tech scmos
magscale 1 2
timestamp 1646624542
<< checkpaint >>
rect -78 -66 116 270
<< nwell >>
rect -18 96 56 210
<< ntransistor >>
rect 14 12 18 52
rect 30 12 34 52
<< ptransistor >>
rect 14 108 18 188
rect 30 108 34 188
<< ndiffusion >>
rect 4 51 14 52
rect 12 13 14 51
rect 4 12 14 13
rect 18 51 30 52
rect 18 13 20 51
rect 28 13 30 51
rect 18 12 30 13
rect 34 51 44 52
rect 34 13 36 51
rect 34 12 44 13
<< pdiffusion >>
rect 4 187 14 188
rect 12 109 14 187
rect 4 108 14 109
rect 18 187 30 188
rect 18 109 20 187
rect 28 109 30 187
rect 18 108 30 109
rect 34 187 44 188
rect 34 109 36 187
rect 34 108 44 109
<< ndcontact >>
rect 4 13 12 51
rect 20 13 28 51
rect 36 13 44 51
<< pdcontact >>
rect 4 109 12 187
rect 20 109 28 187
rect 36 109 44 187
<< psubstratepcontact >>
rect -4 -4 4 4
rect 28 -4 36 4
<< nsubstratencontact >>
rect -4 196 4 204
rect 28 196 36 204
<< polysilicon >>
rect 14 188 18 192
rect 30 188 34 192
rect 14 106 18 108
rect 30 106 34 108
rect 14 102 34 106
rect 14 66 18 102
rect 12 60 18 66
rect 12 58 34 60
rect 14 56 34 58
rect 14 52 18 56
rect 30 52 34 56
rect 14 8 18 12
rect 30 8 34 12
<< polycontact >>
rect 4 58 12 66
<< metal1 >>
rect -4 204 52 206
rect 4 196 28 204
rect 36 196 52 204
rect -4 194 52 196
rect 4 187 12 194
rect 4 108 12 109
rect 20 187 28 188
rect 4 66 12 74
rect 4 51 12 52
rect 4 6 12 13
rect 20 51 28 109
rect 36 187 44 194
rect 36 108 44 109
rect 20 12 28 13
rect 36 51 44 52
rect 36 6 44 13
rect -4 4 52 6
rect 4 -4 28 4
rect 36 -4 52 4
rect -4 -6 52 -4
<< m1p >>
rect 20 86 28 94
rect 4 66 12 74
<< labels >>
rlabel metal1 8 200 8 200 4 vdd
rlabel metal1 8 0 8 0 4 gnd
rlabel metal1 24 90 24 90 4 Y
rlabel metal1 8 70 8 70 4 A
<< end >>
