* NGSPICE file created from address_gen.ext - technology: scmos

* Black-box entry subcircuit for FILL abstract view
.subckt FILL gnd vdd
.ends

* Black-box entry subcircuit for AND2X2 abstract view
.subckt AND2X2 A B gnd Y vdd
.ends

* Black-box entry subcircuit for NAND2X1 abstract view
.subckt NAND2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for OAI21X1 abstract view
.subckt OAI21X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for INVX1 abstract view
.subckt INVX1 A gnd Y vdd
.ends

* Black-box entry subcircuit for OR2X2 abstract view
.subckt OR2X2 A B gnd Y vdd
.ends

* Black-box entry subcircuit for NOR3X1 abstract view
.subckt NOR3X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for CLKBUF1 abstract view
.subckt CLKBUF1 A gnd Y vdd
.ends

* Black-box entry subcircuit for NAND3X1 abstract view
.subckt NAND3X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for DFFPOSX1 abstract view
.subckt DFFPOSX1 Q CLK D gnd vdd
.ends

* Black-box entry subcircuit for BUFX2 abstract view
.subckt BUFX2 A gnd Y vdd
.ends

* Black-box entry subcircuit for AOI21X1 abstract view
.subckt AOI21X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for NOR2X1 abstract view
.subckt NOR2X1 A B gnd Y vdd
.ends

.subckt address_gen vdd gnd address_enable clock reset address_a[0] address_a[1] address_a[2]
+ address_a[3] address_a[4] address_a[5] address_a[6] address_a[7] address_a[8] address_a[9]
+ address_a[10] address_a[11] address_a[12] address_a[13] address_a[14] address_a[15]
+ address_b[0] address_b[1] address_b[2] address_b[3] address_b[4] address_b[5] address_b[6]
+ address_b[7] address_b[8] address_b[9] address_b[10] address_b[11] address_b[12]
+ address_b[13] address_b[14] address_b[15]
XFILL_5_1_2 gnd vdd FILL
XAND2X2_5 BUFX2_24/A BUFX2_25/A gnd AND2X2_5/Y vdd AND2X2
XNAND2X1_10 BUFX2_10/A BUFX2_11/A gnd OAI21X1_7/A vdd NAND2X1
XNAND2X1_21 BUFX2_3/Y NOR3X1_1/C gnd NOR2X1_22/A vdd NAND2X1
XOAI21X1_19 NOR3X1_1/A NOR3X1_1/C OAI21X1_19/C gnd NOR2X1_23/B vdd OAI21X1
XFILL_8_1_0 gnd vdd FILL
XINVX1_6 INVX1_6/A gnd INVX1_6/Y vdd INVX1
XFILL_0_0_0 gnd vdd FILL
XOR2X2_4 OR2X2_4/A OR2X2_4/B gnd OR2X2_4/Y vdd OR2X2
XNAND2X1_11 BUFX2_12/A BUFX2_13/A gnd NOR2X1_11/B vdd NAND2X1
XAND2X2_6 BUFX2_2/Y BUFX2_6/A gnd AND2X2_6/Y vdd AND2X2
XNAND2X1_22 NOR2X1_2/Y NOR2X1_3/Y gnd OAI21X1_22/B vdd NAND2X1
XFILL_0_0_1 gnd vdd FILL
XFILL_8_1_1 gnd vdd FILL
XINVX1_7 INVX1_7/A gnd INVX1_7/Y vdd INVX1
XAND2X2_7 address_enable BUFX2_7/A gnd NOR2X1_5/A vdd AND2X2
XNAND2X1_12 INVX1_7/Y NOR2X1_11/Y gnd OAI21X1_9/B vdd NAND2X1
XFILL_8_1_2 gnd vdd FILL
XINVX1_8 INVX1_8/A gnd INVX1_8/Y vdd INVX1
XFILL_0_0_2 gnd vdd FILL
XAND2X2_8 OR2X2_1/Y AND2X2_8/B gnd AND2X2_8/Y vdd AND2X2
XNAND2X1_13 BUFX2_14/A BUFX2_15/A gnd INVX1_8/A vdd NAND2X1
XNOR3X1_1 NOR3X1_1/A NOR3X1_1/B NOR3X1_1/C gnd NOR3X1_1/Y vdd NOR3X1
XFILL_3_0_0 gnd vdd FILL
XAND2X2_9 OR2X2_2/Y AND2X2_9/B gnd AND2X2_9/Y vdd AND2X2
XINVX1_9 INVX1_9/A gnd OR2X2_1/B vdd INVX1
XNAND2X1_14 BUFX2_5/Y OR2X2_1/A gnd NOR2X1_14/A vdd NAND2X1
XNOR3X1_2 NOR3X1_2/A NOR3X1_2/B NOR3X1_2/C gnd NOR3X1_3/B vdd NOR3X1
XCLKBUF1_1 clock gnd CLKBUF1_1/Y vdd CLKBUF1
XFILL_3_0_1 gnd vdd FILL
XNAND2X1_15 INVX1_9/A INVX1_10/A gnd NOR2X1_15/B vdd NAND2X1
XNOR3X1_3 reset NOR3X1_3/B NOR3X1_3/C gnd NOR3X1_3/Y vdd NOR3X1
XFILL_3_0_2 gnd vdd FILL
XCLKBUF1_2 clock gnd CLKBUF1_2/Y vdd CLKBUF1
XNAND2X1_16 BUFX2_5/Y OR2X2_2/A gnd NAND2X1_16/Y vdd NAND2X1
XNAND3X1_1 AND2X2_3/Y AND2X2_4/Y AND2X2_5/Y gnd NOR3X1_1/C vdd NAND3X1
XFILL_1_1_0 gnd vdd FILL
XFILL_6_0_0 gnd vdd FILL
XCLKBUF1_3 clock gnd CLKBUF1_3/Y vdd CLKBUF1
XNAND3X1_2 INVX1_21/A INVX1_20/A NOR3X1_1/Y gnd NAND3X1_2/Y vdd NAND3X1
XNAND2X1_17 INVX1_11/A INVX1_12/A gnd NOR2X1_18/A vdd NAND2X1
XFILL_1_1_1 gnd vdd FILL
XCLKBUF1_4 clock gnd CLKBUF1_4/Y vdd CLKBUF1
XFILL_6_0_1 gnd vdd FILL
XNAND2X1_18 address_enable BUFX2_20/A gnd NOR2X1_18/B vdd NAND2X1
XFILL_1_1_2 gnd vdd FILL
XNAND3X1_3 NOR2X1_1/Y NOR2X1_2/Y NOR2X1_3/Y gnd NOR3X1_2/C vdd NAND3X1
XFILL_6_0_2 gnd vdd FILL
XCLKBUF1_5 clock gnd CLKBUF1_5/Y vdd CLKBUF1
XFILL_4_1_0 gnd vdd FILL
XNAND3X1_4 INVX1_21/A INVX1_20/A INVX1_1/A gnd NOR2X1_4/A vdd NAND3X1
XOAI21X1_1 NOR2X1_4/A NOR3X1_2/C BUFX2_1/Y gnd OAI21X1_1/Y vdd OAI21X1
XNAND2X1_19 AND2X2_10/Y AND2X2_11/Y gnd OAI21X1_12/B vdd NAND2X1
XFILL_5_1 gnd vdd FILL
XFILL_4_1_1 gnd vdd FILL
XNAND3X1_5 BUFX2_7/A BUFX2_8/A BUFX2_9/A gnd INVX1_7/A vdd NAND3X1
XOAI21X1_2 NOR2X1_4/A NOR3X1_2/C INVX1_3/Y gnd OAI21X1_2/Y vdd OAI21X1
XFILL_4_1_2 gnd vdd FILL
XNAND3X1_6 NOR2X1_11/Y INVX1_8/Y INVX1_6/A gnd OR2X2_1/A vdd NAND3X1
XOAI21X1_3 address_enable BUFX2_7/A BUFX2_3/Y gnd NOR2X1_5/B vdd OAI21X1
XFILL_7_1_0 gnd vdd FILL
XDFFPOSX1_30 INVX1_21/A CLKBUF1_1/Y NOR3X1_3/Y gnd vdd DFFPOSX1
XNAND3X1_7 NOR2X1_11/Y NOR2X1_15/Y INVX1_6/A gnd OR2X2_2/A vdd NAND3X1
XBUFX2_1 INVX1_2/Y gnd BUFX2_1/Y vdd BUFX2
XAOI21X1_1 NAND3X1_2/Y INVX1_1/Y OAI21X1_1/Y gnd AOI21X1_1/Y vdd AOI21X1
XOAI21X1_4 BUFX2_8/A NOR2X1_5/A BUFX2_2/Y gnd NOR2X1_6/A vdd OAI21X1
XBUFX2_30 INVX1_16/A gnd address_b[8] vdd BUFX2
XAOI21X1_20 OR2X2_4/A OR2X2_4/B reset gnd AND2X2_14/B vdd AOI21X1
XDFFPOSX1_31 INVX1_1/A CLKBUF1_1/Y AOI21X1_1/Y gnd vdd DFFPOSX1
XDFFPOSX1_20 BUFX2_25/A CLKBUF1_3/Y NOR2X1_21/Y gnd vdd DFFPOSX1
XFILL_7_1_1 gnd vdd FILL
XAOI21X1_2 INVX1_3/A NOR2X1_4/Y NAND2X1_8/Y gnd AOI21X1_2/Y vdd AOI21X1
XBUFX2_2 INVX1_2/Y gnd BUFX2_2/Y vdd BUFX2
XBUFX2_20 BUFX2_20/A gnd address_a[14] vdd BUFX2
XBUFX2_31 INVX1_17/A gnd address_b[9] vdd BUFX2
XNAND3X1_8 AND2X2_1/Y NOR2X1_2/Y NOR2X1_3/Y gnd OR2X2_4/A vdd NAND3X1
XAOI21X1_10 OR2X2_1/Y INVX1_10/Y NAND2X1_16/Y gnd AOI21X1_10/Y vdd AOI21X1
XOAI21X1_5 BUFX2_9/A INVX1_4/Y BUFX2_2/Y gnd NOR2X1_8/B vdd OAI21X1
XAOI21X1_21 OR2X2_4/Y INVX1_19/Y OAI21X1_22/Y gnd AOI21X1_21/Y vdd AOI21X1
XDFFPOSX1_32 INVX1_3/A CLKBUF1_5/Y AOI21X1_2/Y gnd vdd DFFPOSX1
XFILL_7_1_2 gnd vdd FILL
XDFFPOSX1_10 BUFX2_15/A CLKBUF1_1/Y NOR2X1_14/Y gnd vdd DFFPOSX1
XDFFPOSX1_21 BUFX2_26/A CLKBUF1_2/Y AOI21X1_16/Y gnd vdd DFFPOSX1
XBUFX2_3 INVX1_2/Y gnd BUFX2_3/Y vdd BUFX2
XBUFX2_10 BUFX2_10/A gnd address_a[4] vdd BUFX2
XBUFX2_21 INVX1_13/A gnd address_a[15] vdd BUFX2
XOAI21X1_6 BUFX2_10/A INVX1_6/A BUFX2_1/Y gnd OAI21X1_6/Y vdd OAI21X1
XAOI21X1_3 BUFX2_10/A INVX1_6/A OAI21X1_6/Y gnd AOI21X1_3/Y vdd AOI21X1
XAOI21X1_11 OR2X2_2/A OR2X2_2/B reset gnd AND2X2_9/B vdd AOI21X1
XAOI21X1_22 NOR3X1_2/B NOR3X1_2/C OAI21X1_23/Y gnd AOI21X1_22/Y vdd AOI21X1
XNOR2X1_1 NOR2X1_1/A NOR2X1_1/B gnd NOR2X1_1/Y vdd NOR2X1
XBUFX2_32 INVX1_18/A gnd address_b[10] vdd BUFX2
XDFFPOSX1_11 INVX1_9/A CLKBUF1_4/Y AND2X2_8/Y gnd vdd DFFPOSX1
XFILL_2_0_0 gnd vdd FILL
XDFFPOSX1_22 BUFX2_27/A CLKBUF1_3/Y NOR2X1_22/Y gnd vdd DFFPOSX1
XBUFX2_22 OR2X2_3/B gnd address_b[0] vdd BUFX2
XBUFX2_11 BUFX2_11/A gnd address_a[5] vdd BUFX2
XAOI21X1_4 INVX1_6/A BUFX2_10/A BUFX2_11/A gnd NOR2X1_9/A vdd AOI21X1
XBUFX2_4 INVX1_2/Y gnd BUFX2_4/Y vdd BUFX2
XNOR2X1_2 NOR2X1_2/A NOR3X1_1/A gnd NOR2X1_2/Y vdd NOR2X1
XBUFX2_33 INVX1_19/A gnd address_b[11] vdd BUFX2
XOAI21X1_7 OAI21X1_7/A INVX1_6/Y BUFX2_1/Y gnd NOR2X1_9/B vdd OAI21X1
XAOI21X1_12 OR2X2_2/Y INVX1_12/Y OAI21X1_11/Y gnd AOI21X1_12/Y vdd AOI21X1
XAOI21X1_23 NOR3X1_1/Y INVX1_20/A INVX1_21/A gnd NOR3X1_3/C vdd AOI21X1
XDFFPOSX1_12 INVX1_10/A CLKBUF1_4/Y AOI21X1_10/Y gnd vdd DFFPOSX1
XDFFPOSX1_23 INVX1_14/A CLKBUF1_2/Y AOI21X1_18/Y gnd vdd DFFPOSX1
XFILL_1_1 gnd vdd FILL
XFILL_2_0_1 gnd vdd FILL
XBUFX2_12 BUFX2_12/A gnd address_a[6] vdd BUFX2
XOAI21X1_8 BUFX2_12/A OAI21X1_8/B BUFX2_1/Y gnd OAI21X1_8/Y vdd OAI21X1
XAOI21X1_5 BUFX2_12/A OAI21X1_8/B OAI21X1_8/Y gnd AOI21X1_5/Y vdd AOI21X1
XAOI21X1_13 INVX1_13/Y OAI21X1_12/B OAI21X1_12/Y gnd AOI21X1_13/Y vdd AOI21X1
XBUFX2_34 INVX1_20/A gnd address_b[12] vdd BUFX2
XBUFX2_5 INVX1_2/Y gnd BUFX2_5/Y vdd BUFX2
XBUFX2_23 BUFX2_23/A gnd address_b[1] vdd BUFX2
XNOR2X1_3 NOR2X1_3/A NOR2X1_3/B gnd NOR2X1_3/Y vdd NOR2X1
XDFFPOSX1_13 INVX1_11/A CLKBUF1_5/Y AND2X2_9/Y gnd vdd DFFPOSX1
XDFFPOSX1_24 INVX1_15/A CLKBUF1_2/Y NOR2X1_23/Y gnd vdd DFFPOSX1
XFILL_2_0_2 gnd vdd FILL
XBUFX2_13 BUFX2_13/A gnd address_a[7] vdd BUFX2
XAOI21X1_6 OAI21X1_8/B BUFX2_12/A BUFX2_13/A gnd NOR2X1_12/B vdd AOI21X1
XDFFPOSX1_1 BUFX2_6/A CLKBUF1_4/Y AND2X2_6/Y gnd vdd DFFPOSX1
XBUFX2_6 BUFX2_6/A gnd address_a[0] vdd BUFX2
XBUFX2_35 INVX1_21/A gnd address_b[13] vdd BUFX2
XBUFX2_24 BUFX2_24/A gnd address_b[2] vdd BUFX2
XFILL_0_1_0 gnd vdd FILL
XNAND2X1_1 AND2X2_1/Y AND2X2_2/Y gnd NOR3X1_1/B vdd NAND2X1
XNOR2X1_4 NOR2X1_4/A NOR3X1_2/C gnd NOR2X1_4/Y vdd NOR2X1
XOAI21X1_9 INVX1_5/Y OAI21X1_9/B BUFX2_2/Y gnd OAI21X1_9/Y vdd OAI21X1
XAOI21X1_14 BUFX2_24/A AND2X2_4/Y OAI21X1_14/Y gnd AOI21X1_14/Y vdd AOI21X1
XDFFPOSX1_14 INVX1_12/A CLKBUF1_4/Y AOI21X1_12/Y gnd vdd DFFPOSX1
XFILL_5_0_0 gnd vdd FILL
XDFFPOSX1_25 INVX1_16/A CLKBUF1_1/Y AOI21X1_19/Y gnd vdd DFFPOSX1
XAOI21X1_7 BUFX2_14/A NOR2X1_13/Y AOI21X1_7/C gnd AOI21X1_7/Y vdd AOI21X1
XBUFX2_14 BUFX2_14/A gnd address_a[8] vdd BUFX2
XBUFX2_36 INVX1_1/A gnd address_b[14] vdd BUFX2
XAOI21X1_15 AND2X2_4/Y BUFX2_24/A BUFX2_25/A gnd NOR2X1_21/B vdd AOI21X1
XBUFX2_25 BUFX2_25/A gnd address_b[3] vdd BUFX2
XNAND2X1_2 INVX1_15/A INVX1_14/A gnd NOR3X1_1/A vdd NAND2X1
XFILL_0_1_1 gnd vdd FILL
XBUFX2_7 BUFX2_7/A gnd address_a[1] vdd BUFX2
XDFFPOSX1_2 BUFX2_7/A CLKBUF1_3/Y NOR2X1_5/Y gnd vdd DFFPOSX1
XNOR2X1_5 NOR2X1_5/A NOR2X1_5/B gnd NOR2X1_5/Y vdd NOR2X1
XFILL_5_0_1 gnd vdd FILL
XDFFPOSX1_15 BUFX2_20/A CLKBUF1_1/Y NOR2X1_19/Y gnd vdd DFFPOSX1
XDFFPOSX1_26 INVX1_17/A CLKBUF1_2/Y AND2X2_13/Y gnd vdd DFFPOSX1
XAOI21X1_8 NOR2X1_13/Y BUFX2_14/A BUFX2_15/A gnd NOR2X1_14/B vdd AOI21X1
XNAND2X1_3 INVX1_17/A INVX1_16/A gnd NOR2X1_1/A vdd NAND2X1
XFILL_0_1_2 gnd vdd FILL
XBUFX2_8 BUFX2_8/A gnd address_a[2] vdd BUFX2
XBUFX2_15 BUFX2_15/A gnd address_a[9] vdd BUFX2
XBUFX2_37 INVX1_3/A gnd address_b[15] vdd BUFX2
XDFFPOSX1_3 BUFX2_8/A CLKBUF1_3/Y NOR2X1_6/Y gnd vdd DFFPOSX1
XNOR2X1_6 NOR2X1_6/A INVX1_4/Y gnd NOR2X1_6/Y vdd NOR2X1
XBUFX2_26 BUFX2_26/A gnd address_b[4] vdd BUFX2
XAOI21X1_16 BUFX2_26/A NOR2X1_3/Y OAI21X1_16/Y gnd AOI21X1_16/Y vdd AOI21X1
XDFFPOSX1_16 INVX1_13/A CLKBUF1_1/Y AOI21X1_13/Y gnd vdd DFFPOSX1
XFILL_5_0_2 gnd vdd FILL
XDFFPOSX1_27 INVX1_18/A CLKBUF1_2/Y AND2X2_14/Y gnd vdd DFFPOSX1
XFILL_3_1_0 gnd vdd FILL
XBUFX2_16 INVX1_9/A gnd address_a[10] vdd BUFX2
XAOI21X1_9 OR2X2_1/A OR2X2_1/B reset gnd AND2X2_8/B vdd AOI21X1
XNOR2X1_7 INVX1_5/Y INVX1_7/A gnd INVX1_6/A vdd NOR2X1
XDFFPOSX1_4 BUFX2_9/A CLKBUF1_4/Y NOR2X1_8/Y gnd vdd DFFPOSX1
XBUFX2_9 BUFX2_9/A gnd address_a[3] vdd BUFX2
XBUFX2_27 BUFX2_27/A gnd address_b[5] vdd BUFX2
XAOI21X1_17 NOR2X1_3/Y BUFX2_26/A BUFX2_27/A gnd NOR2X1_22/B vdd AOI21X1
XNAND2X1_4 INVX1_19/A INVX1_18/A gnd NOR2X1_1/B vdd NAND2X1
XFILL_8_0_0 gnd vdd FILL
XDFFPOSX1_17 OR2X2_3/B CLKBUF1_5/Y OR2X2_3/Y gnd vdd DFFPOSX1
XDFFPOSX1_28 INVX1_19/A CLKBUF1_2/Y AOI21X1_21/Y gnd vdd DFFPOSX1
XFILL_3_1_1 gnd vdd FILL
XNAND2X1_5 BUFX2_27/A BUFX2_26/A gnd NOR2X1_2/A vdd NAND2X1
XDFFPOSX1_5 BUFX2_10/A CLKBUF1_5/Y AOI21X1_3/Y gnd vdd DFFPOSX1
XFILL_8_0_1 gnd vdd FILL
XBUFX2_17 INVX1_10/A gnd address_a[11] vdd BUFX2
XINVX1_20 INVX1_20/A gnd NOR3X1_2/B vdd INVX1
XNOR2X1_8 INVX1_6/A NOR2X1_8/B gnd NOR2X1_8/Y vdd NOR2X1
XAOI21X1_18 INVX1_14/Y NOR3X1_1/C OAI21X1_17/Y gnd AOI21X1_18/Y vdd AOI21X1
XBUFX2_28 INVX1_14/A gnd address_b[6] vdd BUFX2
XDFFPOSX1_29 INVX1_20/A CLKBUF1_2/Y AOI21X1_22/Y gnd vdd DFFPOSX1
XDFFPOSX1_18 BUFX2_23/A CLKBUF1_3/Y NOR2X1_20/Y gnd vdd DFFPOSX1
XBUFX2_18 INVX1_11/A gnd address_a[12] vdd BUFX2
XDFFPOSX1_6 BUFX2_11/A CLKBUF1_5/Y NOR2X1_9/Y gnd vdd DFFPOSX1
XNOR2X1_9 NOR2X1_9/A NOR2X1_9/B gnd NOR2X1_9/Y vdd NOR2X1
XINVX1_10 INVX1_10/A gnd INVX1_10/Y vdd INVX1
XINVX1_21 INVX1_21/A gnd NOR3X1_2/A vdd INVX1
XFILL_3_1_2 gnd vdd FILL
XNAND2X1_6 BUFX2_23/A address_enable gnd NOR2X1_3/A vdd NAND2X1
XBUFX2_29 INVX1_15/A gnd address_b[7] vdd BUFX2
XFILL_8_0_2 gnd vdd FILL
XAOI21X1_19 INVX1_16/Y OAI21X1_22/B OAI21X1_20/Y gnd AOI21X1_19/Y vdd AOI21X1
XDFFPOSX1_19 BUFX2_24/A CLKBUF1_3/Y AOI21X1_14/Y gnd vdd DFFPOSX1
XFILL_6_1_0 gnd vdd FILL
XNAND2X1_7 BUFX2_24/A BUFX2_25/A gnd NOR2X1_3/B vdd NAND2X1
XDFFPOSX1_7 BUFX2_12/A CLKBUF1_5/Y AOI21X1_5/Y gnd vdd DFFPOSX1
XBUFX2_19 INVX1_12/A gnd address_a[13] vdd BUFX2
XINVX1_11 INVX1_11/A gnd OR2X2_2/B vdd INVX1
XFILL_6_1_1 gnd vdd FILL
XINVX1_12 INVX1_12/A gnd INVX1_12/Y vdd INVX1
XNAND2X1_8 BUFX2_1/Y OAI21X1_2/Y gnd NAND2X1_8/Y vdd NAND2X1
XDFFPOSX1_8 BUFX2_13/A CLKBUF1_1/Y NOR2X1_12/Y gnd vdd DFFPOSX1
XNOR2X1_20 AND2X2_4/Y NOR2X1_20/B gnd NOR2X1_20/Y vdd NOR2X1
XAND2X2_10 NOR2X1_18/Y INVX1_7/Y gnd AND2X2_10/Y vdd AND2X2
XNOR2X1_10 OAI21X1_7/A INVX1_6/Y gnd OAI21X1_8/B vdd NOR2X1
XFILL_6_1_2 gnd vdd FILL
XNOR2X1_21 NOR2X1_21/A NOR2X1_21/B gnd NOR2X1_21/Y vdd NOR2X1
XDFFPOSX1_9 BUFX2_14/A CLKBUF1_4/Y AOI21X1_7/Y gnd vdd DFFPOSX1
XINVX1_13 INVX1_13/A gnd INVX1_13/Y vdd INVX1
XNAND2X1_9 BUFX2_8/A NOR2X1_5/A gnd INVX1_4/A vdd NAND2X1
XFILL_6_1 gnd vdd FILL
XAND2X2_11 NOR2X1_11/Y NOR2X1_15/Y gnd AND2X2_11/Y vdd AND2X2
XFILL_1_0_0 gnd vdd FILL
XNOR2X1_11 OAI21X1_7/A NOR2X1_11/B gnd NOR2X1_11/Y vdd NOR2X1
XINVX1_14 INVX1_14/A gnd INVX1_14/Y vdd INVX1
XNOR2X1_22 NOR2X1_22/A NOR2X1_22/B gnd NOR2X1_22/Y vdd NOR2X1
XOAI21X1_20 INVX1_16/Y OAI21X1_22/B BUFX2_4/Y gnd OAI21X1_20/Y vdd OAI21X1
XFILL_1_0_1 gnd vdd FILL
XAND2X2_12 OR2X2_4/A BUFX2_4/Y gnd AND2X2_13/A vdd AND2X2
XNOR2X1_12 OAI21X1_9/Y NOR2X1_12/B gnd NOR2X1_12/Y vdd NOR2X1
XINVX1_15 INVX1_15/A gnd INVX1_15/Y vdd INVX1
XNOR2X1_23 reset NOR2X1_23/B gnd NOR2X1_23/Y vdd NOR2X1
XOAI21X1_10 BUFX2_14/A NOR2X1_13/Y BUFX2_2/Y gnd AOI21X1_7/C vdd OAI21X1
XAND2X2_13 AND2X2_13/A AND2X2_13/B gnd AND2X2_13/Y vdd AND2X2
XOAI21X1_21 INVX1_16/Y OAI21X1_22/B INVX1_17/Y gnd AND2X2_13/B vdd OAI21X1
XFILL_1_0_2 gnd vdd FILL
XNOR2X1_13 INVX1_5/Y OAI21X1_9/B gnd NOR2X1_13/Y vdd NOR2X1
XINVX1_16 INVX1_16/A gnd INVX1_16/Y vdd INVX1
XOAI21X1_11 NOR2X1_18/A OR2X2_2/A BUFX2_5/Y gnd OAI21X1_11/Y vdd OAI21X1
XOAI21X1_22 NOR3X1_1/B OAI21X1_22/B BUFX2_4/Y gnd OAI21X1_22/Y vdd OAI21X1
XFILL_4_0_0 gnd vdd FILL
XAND2X2_14 OR2X2_4/Y AND2X2_14/B gnd AND2X2_14/Y vdd AND2X2
XFILL_4_1 gnd vdd FILL
XNOR2X1_14 NOR2X1_14/A NOR2X1_14/B gnd NOR2X1_14/Y vdd NOR2X1
XINVX1_17 INVX1_17/A gnd INVX1_17/Y vdd INVX1
XOAI21X1_12 INVX1_13/Y OAI21X1_12/B BUFX2_5/Y gnd OAI21X1_12/Y vdd OAI21X1
XOAI21X1_23 NOR3X1_2/B NOR3X1_2/C BUFX2_1/Y gnd OAI21X1_23/Y vdd OAI21X1
XFILL_4_0_1 gnd vdd FILL
XNOR2X1_15 INVX1_8/A NOR2X1_15/B gnd NOR2X1_15/Y vdd NOR2X1
XINVX1_18 INVX1_18/A gnd OR2X2_4/B vdd INVX1
XFILL_4_0_2 gnd vdd FILL
XOAI21X1_13 BUFX2_23/A address_enable BUFX2_3/Y gnd NOR2X1_20/B vdd OAI21X1
XNOR2X1_16 NOR2X1_18/A OR2X2_2/A gnd NOR2X1_17/B vdd NOR2X1
XINVX1_19 INVX1_19/A gnd INVX1_19/Y vdd INVX1
XFILL_2_1_0 gnd vdd FILL
XFILL_7_0_0 gnd vdd FILL
XOAI21X1_14 BUFX2_24/A AND2X2_4/Y BUFX2_3/Y gnd OAI21X1_14/Y vdd OAI21X1
XINVX1_1 INVX1_1/A gnd INVX1_1/Y vdd INVX1
XNOR2X1_17 BUFX2_20/A NOR2X1_17/B gnd NOR2X1_19/B vdd NOR2X1
XFILL_2_1 gnd vdd FILL
XFILL_2_1_1 gnd vdd FILL
XAND2X2_1 INVX1_17/A INVX1_16/A gnd AND2X2_1/Y vdd AND2X2
XFILL_7_0_1 gnd vdd FILL
XOAI21X1_15 NOR2X1_3/A NOR2X1_3/B BUFX2_3/Y gnd NOR2X1_21/A vdd OAI21X1
XINVX1_2 reset gnd INVX1_2/Y vdd INVX1
XAND2X2_2 INVX1_19/A INVX1_18/A gnd AND2X2_2/Y vdd AND2X2
XNOR2X1_18 NOR2X1_18/A NOR2X1_18/B gnd NOR2X1_18/Y vdd NOR2X1
XFILL_2_2 gnd vdd FILL
XFILL_2_1_2 gnd vdd FILL
XFILL_7_0_2 gnd vdd FILL
XOAI21X1_16 BUFX2_26/A NOR2X1_3/Y BUFX2_4/Y gnd OAI21X1_16/Y vdd OAI21X1
XOR2X2_1 OR2X2_1/A OR2X2_1/B gnd OR2X2_1/Y vdd OR2X2
XINVX1_3 INVX1_3/A gnd INVX1_3/Y vdd INVX1
XFILL_5_1_0 gnd vdd FILL
XNOR2X1_19 NOR2X1_19/A NOR2X1_19/B gnd NOR2X1_19/Y vdd NOR2X1
XAND2X2_3 BUFX2_27/A BUFX2_26/A gnd AND2X2_3/Y vdd AND2X2
XOAI21X1_17 INVX1_14/Y NOR3X1_1/C BUFX2_4/Y gnd OAI21X1_17/Y vdd OAI21X1
XOR2X2_2 OR2X2_2/A OR2X2_2/B gnd OR2X2_2/Y vdd OR2X2
XFILL_5_1_1 gnd vdd FILL
XINVX1_4 INVX1_4/A gnd INVX1_4/Y vdd INVX1
XNAND2X1_20 BUFX2_5/Y OAI21X1_12/B gnd NOR2X1_19/A vdd NAND2X1
XAND2X2_4 BUFX2_23/A address_enable gnd AND2X2_4/Y vdd AND2X2
XOAI21X1_18 INVX1_14/Y NOR3X1_1/C INVX1_15/Y gnd OAI21X1_19/C vdd OAI21X1
XOR2X2_3 reset OR2X2_3/B gnd OR2X2_3/Y vdd OR2X2
XINVX1_5 address_enable gnd INVX1_5/Y vdd INVX1
.ends

