* NGSPICE file created from sigmoid_approx.ext - technology: scmos

* Black-box entry subcircuit for FILL abstract view
.subckt FILL gnd vdd
.ends

* Black-box entry subcircuit for AND2X2 abstract view
.subckt AND2X2 A B gnd Y vdd
.ends

* Black-box entry subcircuit for NAND2X1 abstract view
.subckt NAND2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for XNOR2X1 abstract view
.subckt XNOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for INVX1 abstract view
.subckt INVX1 A gnd Y vdd
.ends

* Black-box entry subcircuit for AOI22X1 abstract view
.subckt AOI22X1 A B C D gnd Y vdd
.ends

* Black-box entry subcircuit for NOR3X1 abstract view
.subckt NOR3X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for MUX2X1 abstract view
.subckt MUX2X1 A B S gnd Y vdd
.ends

* Black-box entry subcircuit for NAND3X1 abstract view
.subckt NAND3X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for XOR2X1 abstract view
.subckt XOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for OAI21X1 abstract view
.subckt OAI21X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for BUFX2 abstract view
.subckt BUFX2 A gnd Y vdd
.ends

* Black-box entry subcircuit for AOI21X1 abstract view
.subckt AOI21X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for NOR2X1 abstract view
.subckt NOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for OR2X2 abstract view
.subckt OR2X2 A B gnd Y vdd
.ends

* Black-box entry subcircuit for OAI22X1 abstract view
.subckt OAI22X1 A B C D gnd Y vdd
.ends

.subckt sigmoid_approx vdd gnd Y[0] Y[1] Y[2] Y[3] Y[4] Y[5] Y[6] Y[7] Y[8] Y[9] Y[10]
+ Y[11] Y[12] Y[13] Y[14] Y[15] Y[16] Y[17] Y[18] Y[19] Y[20] Y[21] Y[22] Y[23] Y[24]
+ Y[25] Y[26] Y[27] Y[28] Y[29] Y[30] Y[31] O[0] O[1] O[2] O[3] O[4] O[5] O[6] O[7]
+ O[8] O[9] O[10] O[11] O[12] O[13] O[14] O[15] O[16] O[17] O[18] O[19] O[20] O[21]
+ O[22] O[23] O[24] O[25] O[26] O[27] O[28] O[29] O[30] O[31]
XFILL_5_1_2 gnd vdd FILL
XAND2X2_5 AND2X2_5/A AND2X2_5/B gnd AND2X2_5/Y vdd AND2X2
XNAND2X1_10 AND2X2_3/Y AND2X2_4/Y gnd NOR3X1_2/B vdd NAND2X1
XXNOR2X1_6 XNOR2X1_6/A Y[9] gnd NOR3X1_9/B vdd XNOR2X1
XINVX1_6 Y[26] gnd INVX1_6/Y vdd INVX1
XFILL_0_0_0 gnd vdd FILL
XAOI22X1_1 OR2X2_2/A OAI21X1_2/Y AOI22X1_1/C OAI21X1_3/Y gnd AOI22X1_1/Y vdd AOI22X1
XAND2X2_6 INVX1_4/A AND2X2_6/B gnd AND2X2_6/Y vdd AND2X2
XNAND2X1_11 AND2X2_5/Y AND2X2_6/Y gnd NOR3X1_2/C vdd NAND2X1
XFILL_0_0_1 gnd vdd FILL
XXNOR2X1_7 XNOR2X1_7/A INVX1_12/Y gnd XNOR2X1_7/Y vdd XNOR2X1
XINVX1_7 Y[28] gnd INVX1_7/Y vdd INVX1
XAND2X2_7 OR2X2_2/Y AND2X2_7/B gnd AND2X2_7/Y vdd AND2X2
XNAND2X1_12 INVX1_3/A NOR3X1_2/Y gnd AOI22X1_1/C vdd NAND2X1
XAOI22X1_2 INVX1_14/A OAI21X1_5/Y BUFX2_6/Y OAI22X1_1/Y gnd AOI22X1_2/Y vdd AOI22X1
XINVX1_8 Y[18] gnd INVX1_8/Y vdd INVX1
XFILL_0_0_2 gnd vdd FILL
XXNOR2X1_8 XNOR2X1_8/A Y[15] gnd XNOR2X1_8/Y vdd XNOR2X1
XAND2X2_8 Y[21] Y[22] gnd MUX2X1_1/A vdd AND2X2
XNOR3X1_1 Y[28] INVX1_3/Y OR2X2_2/A gnd NOR3X1_1/Y vdd NOR3X1
XNAND2X1_13 Y[18] OAI21X1_4/Y gnd NAND2X1_14/B vdd NAND2X1
XFILL_3_0_0 gnd vdd FILL
XAND2X2_9 AND2X2_9/A AND2X2_9/B gnd AND2X2_9/Y vdd AND2X2
XINVX1_9 Y[16] gnd INVX1_9/Y vdd INVX1
XNOR3X1_2 NOR3X1_2/A NOR3X1_2/B NOR3X1_2/C gnd NOR3X1_2/Y vdd NOR3X1
XNAND2X1_14 NAND3X1_4/Y NAND2X1_14/B gnd INVX1_14/A vdd NAND2X1
XFILL_3_0_1 gnd vdd FILL
XNOR3X1_3 Y[26] OR2X2_2/B OR2X2_2/A gnd NOR3X1_3/Y vdd NOR3X1
XNAND2X1_15 BUFX2_7/Y NOR2X1_5/A gnd XOR2X1_1/A vdd NAND2X1
XMUX2X1_1 MUX2X1_1/A INVX1_4/A MUX2X1_1/S gnd MUX2X1_1/Y vdd MUX2X1
XFILL_3_0_2 gnd vdd FILL
XNOR3X1_4 NOR3X1_9/A XOR2X1_1/Y BUFX2_2/Y gnd BUFX2_9/A vdd NOR3X1
XNAND2X1_16 NOR2X1_3/Y AND2X2_1/Y gnd OAI21X1_10/B vdd NAND2X1
XNAND3X1_1 NOR2X1_5/Y NOR2X1_10/Y NOR2X1_15/Y gnd OR2X2_2/A vdd NAND3X1
XFILL_1_1_0 gnd vdd FILL
XFILL_6_0_0 gnd vdd FILL
XXOR2X1_1 XOR2X1_1/A Y[4] gnd XOR2X1_1/Y vdd XOR2X1
XNAND3X1_2 INVX1_5/Y AND2X2_5/Y NOR2X1_19/Y gnd MUX2X1_1/S vdd NAND3X1
XNOR3X1_5 NOR3X1_9/A XOR2X1_2/Y BUFX2_2/Y gnd NOR3X1_5/Y vdd NOR3X1
XNAND2X1_17 INVX1_1/A OAI21X1_10/B gnd XOR2X1_3/A vdd NAND2X1
XFILL_1_1_1 gnd vdd FILL
XFILL_6_0_1 gnd vdd FILL
XXOR2X1_2 XOR2X1_2/A Y[5] gnd XOR2X1_2/Y vdd XOR2X1
XNAND3X1_3 AND2X2_5/A NOR2X1_5/Y NOR2X1_10/Y gnd OAI21X1_8/B vdd NAND3X1
XFILL_1_1_2 gnd vdd FILL
XNOR3X1_6 NOR3X1_9/A XOR2X1_3/Y BUFX2_4/Y gnd NOR3X1_6/Y vdd NOR3X1
XNAND2X1_18 NOR2X1_6/Y NOR2X1_5/Y gnd OAI21X1_13/B vdd NAND2X1
XFILL_6_0_2 gnd vdd FILL
XXOR2X1_3 XOR2X1_3/A Y[6] gnd XOR2X1_3/Y vdd XOR2X1
XFILL_4_1_0 gnd vdd FILL
XOAI21X1_1 NOR3X1_1/Y OAI21X1_1/B OAI21X1_1/C gnd OAI21X1_1/Y vdd OAI21X1
XFILL_5_1 gnd vdd FILL
XNAND3X1_4 BUFX2_6/Y INVX1_8/Y OAI21X1_8/B gnd NAND3X1_4/Y vdd NAND3X1
XNAND2X1_19 BUFX2_8/Y OAI21X1_13/B gnd XOR2X1_5/A vdd NAND2X1
XNOR3X1_7 NOR3X1_9/A XOR2X1_4/Y BUFX2_4/Y gnd NOR3X1_7/Y vdd NOR3X1
XXOR2X1_4 XOR2X1_4/A Y[7] gnd XOR2X1_4/Y vdd XOR2X1
XFILL_4_1_1 gnd vdd FILL
XNAND3X1_5 INVX1_9/Y NOR2X1_5/Y NOR2X1_10/Y gnd OAI21X1_4/B vdd NAND3X1
XNOR3X1_8 NOR3X1_9/A NOR3X1_8/B BUFX2_2/Y gnd NOR3X1_8/Y vdd NOR3X1
XOAI21X1_2 INVX1_4/Y MUX2X1_1/S Y[23] gnd OAI21X1_2/Y vdd OAI21X1
XXOR2X1_5 XOR2X1_5/A Y[10] gnd XOR2X1_5/Y vdd XOR2X1
XFILL_4_1_2 gnd vdd FILL
XBUFX2_40 gnd gnd O[31] vdd BUFX2
XNOR3X1_9 NOR3X1_9/A NOR3X1_9/B BUFX2_2/Y gnd NOR3X1_9/Y vdd NOR3X1
XNAND3X1_6 BUFX2_8/Y Y[17] OAI21X1_4/B gnd INVX1_10/A vdd NAND3X1
XOAI21X1_3 Y[26] OR2X2_2/Y Y[27] gnd OAI21X1_3/Y vdd OAI21X1
XXOR2X1_6 XOR2X1_6/A Y[11] gnd XOR2X1_6/Y vdd XOR2X1
XNAND3X1_7 AND2X2_6/Y AND2X2_9/Y INVX1_3/A gnd NAND3X1_7/Y vdd NAND3X1
XBUFX2_1 BUFX2_4/A gnd BUFX2_1/Y vdd BUFX2
XAOI21X1_1 AOI22X1_1/Y OAI21X1_1/Y INVX1_1/Y gnd NOR3X1_9/A vdd AOI21X1
XBUFX2_30 gnd gnd O[21] vdd BUFX2
XOAI21X1_4 Y[17] OAI21X1_4/B BUFX2_7/Y gnd OAI21X1_4/Y vdd OAI21X1
XFILL_3_1 gnd vdd FILL
XXOR2X1_7 XOR2X1_7/A Y[12] gnd XOR2X1_7/Y vdd XOR2X1
XAOI21X1_2 NOR3X1_2/Y INVX1_2/A INVX1_6/Y gnd OAI22X1_1/B vdd AOI21X1
XBUFX2_2 BUFX2_4/A gnd BUFX2_2/Y vdd BUFX2
XNAND3X1_8 AND2X2_5/Y NOR2X1_5/Y NOR2X1_10/Y gnd XNOR2X1_4/A vdd NAND3X1
XBUFX2_20 BUFX2_20/A gnd O[11] vdd BUFX2
XBUFX2_31 gnd gnd O[22] vdd BUFX2
XOAI21X1_5 OR2X2_3/A OR2X2_3/B XNOR2X1_1/Y gnd OAI21X1_5/Y vdd OAI21X1
XXOR2X1_8 XOR2X1_8/A Y[13] gnd XOR2X1_8/Y vdd XOR2X1
XNAND3X1_9 BUFX2_6/Y XNOR2X1_4/Y XNOR2X1_3/Y gnd NAND3X1_9/Y vdd NAND3X1
XNOR3X1_10 NOR3X1_9/A XOR2X1_5/Y BUFX2_1/Y gnd BUFX2_15/A vdd NOR3X1
XBUFX2_3 BUFX2_4/A gnd BUFX2_3/Y vdd BUFX2
XAOI21X1_3 NOR3X1_2/Y INVX1_3/A INVX1_7/Y gnd OAI22X1_1/D vdd AOI21X1
XOAI21X1_6 Y[24] OR2X2_2/A Y[25] gnd AND2X2_7/B vdd OAI21X1
XNOR2X1_1 Y[0] Y[3] gnd NOR2X1_1/Y vdd NOR2X1
XBUFX2_10 NOR3X1_5/Y gnd O[1] vdd BUFX2
XBUFX2_21 BUFX2_21/A gnd O[12] vdd BUFX2
XBUFX2_32 gnd gnd O[23] vdd BUFX2
XFILL_2_0_0 gnd vdd FILL
XNOR3X1_11 NOR3X1_9/A XOR2X1_6/Y BUFX2_4/Y gnd BUFX2_16/A vdd NOR3X1
XNOR2X1_2 Y[1] Y[2] gnd NOR2X1_2/Y vdd NOR2X1
XBUFX2_33 gnd gnd O[24] vdd BUFX2
XBUFX2_22 BUFX2_22/A gnd O[13] vdd BUFX2
XAOI21X1_4 OAI21X1_4/B INVX1_1/A Y[17] gnd OR2X2_3/B vdd AOI21X1
XBUFX2_11 NOR3X1_6/Y gnd O[2] vdd BUFX2
XBUFX2_4 BUFX2_4/A gnd BUFX2_4/Y vdd BUFX2
XOAI21X1_7 AND2X2_7/Y MUX2X1_1/Y BUFX2_7/Y gnd OAI21X1_7/Y vdd OAI21X1
XFILL_1_1 gnd vdd FILL
XFILL_2_0_1 gnd vdd FILL
XNOR3X1_12 NOR3X1_9/A XOR2X1_7/Y BUFX2_1/Y gnd BUFX2_17/A vdd NOR3X1
XBUFX2_34 gnd gnd O[25] vdd BUFX2
XBUFX2_5 Y[31] gnd INVX1_1/A vdd BUFX2
XOAI21X1_8 Y[18] OAI21X1_8/B BUFX2_8/Y gnd XNOR2X1_2/A vdd OAI21X1
XBUFX2_23 BUFX2_23/A gnd O[14] vdd BUFX2
XAOI21X1_5 NOR2X1_10/Y NOR2X1_5/Y INVX1_1/Y gnd XNOR2X1_1/A vdd AOI21X1
XBUFX2_12 NOR3X1_7/Y gnd O[3] vdd BUFX2
XNOR2X1_3 Y[5] Y[4] gnd NOR2X1_3/Y vdd NOR2X1
XFILL_2_0_2 gnd vdd FILL
XBUFX2_13 NOR3X1_8/Y gnd O[4] vdd BUFX2
XNAND2X1_1 NOR2X1_1/Y NOR2X1_2/Y gnd NOR2X1_5/A vdd NAND2X1
XBUFX2_35 gnd gnd O[26] vdd BUFX2
XBUFX2_6 Y[31] gnd BUFX2_6/Y vdd BUFX2
XAOI21X1_6 NAND3X1_9/Y NAND3X1_7/Y XNOR2X1_2/Y gnd AOI21X1_6/Y vdd AOI21X1
XFILL_0_1_0 gnd vdd FILL
XNOR3X1_13 NOR3X1_9/A XOR2X1_8/Y BUFX2_4/Y gnd BUFX2_18/A vdd NOR3X1
XBUFX2_24 BUFX2_24/A gnd O[15] vdd BUFX2
XOAI21X1_9 Y[4] NOR2X1_5/A BUFX2_8/Y gnd XOR2X1_2/A vdd OAI21X1
XNOR2X1_4 Y[6] Y[7] gnd NOR2X1_4/Y vdd NOR2X1
XFILL_5_0_0 gnd vdd FILL
XNOR3X1_14 NOR3X1_9/A XNOR2X1_7/Y BUFX2_1/Y gnd BUFX2_19/A vdd NOR3X1
XBUFX2_14 NOR3X1_9/Y gnd O[5] vdd BUFX2
XNAND2X1_2 NOR2X1_3/Y NOR2X1_4/Y gnd NOR2X1_5/B vdd NAND2X1
XNOR2X1_5 NOR2X1_5/A NOR2X1_5/B gnd NOR2X1_5/Y vdd NOR2X1
XBUFX2_7 Y[31] gnd BUFX2_7/Y vdd BUFX2
XBUFX2_36 gnd gnd O[27] vdd BUFX2
XBUFX2_25 BUFX2_25/A gnd O[16] vdd BUFX2
XFILL_0_1_1 gnd vdd FILL
XFILL_5_0_1 gnd vdd FILL
XBUFX2_8 Y[31] gnd BUFX2_8/Y vdd BUFX2
XNOR3X1_15 NOR3X1_9/A XNOR2X1_8/Y BUFX2_3/Y gnd BUFX2_20/A vdd NOR3X1
XFILL_0_1_2 gnd vdd FILL
XNAND2X1_3 NOR2X1_6/Y NOR2X1_7/Y gnd NOR2X1_10/A vdd NAND2X1
XBUFX2_37 gnd gnd O[28] vdd BUFX2
XNOR2X1_6 Y[8] Y[9] gnd NOR2X1_6/Y vdd NOR2X1
XBUFX2_26 gnd gnd O[17] vdd BUFX2
XBUFX2_15 BUFX2_15/A gnd O[6] vdd BUFX2
XFILL_5_0_2 gnd vdd FILL
XFILL_3_1_0 gnd vdd FILL
XNOR3X1_16 NOR3X1_9/A XNOR2X1_1/Y BUFX2_3/Y gnd BUFX2_21/A vdd NOR3X1
XBUFX2_38 gnd gnd O[29] vdd BUFX2
XBUFX2_27 gnd gnd O[18] vdd BUFX2
XBUFX2_9 BUFX2_9/A gnd O[0] vdd BUFX2
XNAND2X1_4 NOR2X1_8/Y NOR2X1_9/Y gnd NOR2X1_10/B vdd NAND2X1
XNOR2X1_7 Y[10] Y[11] gnd NOR2X1_7/Y vdd NOR2X1
XBUFX2_16 BUFX2_16/A gnd O[7] vdd BUFX2
XFILL_3_1_1 gnd vdd FILL
XNOR3X1_17 NOR3X1_9/A OR2X2_3/Y BUFX2_3/Y gnd BUFX2_22/A vdd NOR3X1
XNAND2X1_5 AND2X2_5/A AND2X2_5/B gnd NOR2X1_15/A vdd NAND2X1
XBUFX2_39 gnd gnd O[30] vdd BUFX2
XBUFX2_28 gnd gnd O[19] vdd BUFX2
XNOR2X1_8 Y[12] Y[13] gnd NOR2X1_8/Y vdd NOR2X1
XBUFX2_17 BUFX2_17/A gnd O[8] vdd BUFX2
XNOR3X1_18 NOR3X1_9/A INVX1_14/Y BUFX2_1/Y gnd BUFX2_23/A vdd NOR3X1
XNAND2X1_6 INVX1_4/A AND2X2_6/B gnd NOR2X1_15/B vdd NAND2X1
XFILL_3_1_2 gnd vdd FILL
XINVX1_10 INVX1_10/A gnd OR2X2_3/A vdd INVX1
XNOR2X1_9 Y[14] Y[15] gnd NOR2X1_9/Y vdd NOR2X1
XBUFX2_18 BUFX2_18/A gnd O[9] vdd BUFX2
XBUFX2_29 gnd gnd O[20] vdd BUFX2
XFILL_6_1_0 gnd vdd FILL
XNAND2X1_7 Y[30] Y[29] gnd OAI21X1_1/B vdd NAND2X1
XINVX1_11 Y[8] gnd INVX1_11/Y vdd INVX1
XBUFX2_19 BUFX2_19/A gnd O[10] vdd BUFX2
XFILL_6_1_1 gnd vdd FILL
XNOR2X1_20 INVX1_1/A Y[28] gnd AND2X2_9/B vdd NOR2X1
XNAND2X1_8 AND2X2_9/A NOR3X1_1/Y gnd OAI21X1_1/C vdd NAND2X1
XINVX1_12 Y[14] gnd INVX1_12/Y vdd INVX1
XAND2X2_10 BUFX2_3/Y INVX1_1/Y gnd BUFX2_25/A vdd AND2X2
XFILL_6_1_2 gnd vdd FILL
XNAND3X1_10 OAI21X1_7/Y AOI21X1_6/Y AOI22X1_2/Y gnd BUFX2_4/A vdd NAND3X1
XNOR2X1_10 NOR2X1_10/A NOR2X1_10/B gnd NOR2X1_10/Y vdd NOR2X1
XNOR2X1_21 INVX1_1/A BUFX2_1/Y gnd BUFX2_24/A vdd NOR2X1
XNAND2X1_9 AND2X2_1/Y AND2X2_2/Y gnd NOR3X1_2/A vdd NAND2X1
XINVX1_13 NOR2X1_8/Y gnd INVX1_13/Y vdd INVX1
XFILL_6_1 gnd vdd FILL
XFILL_1_0_0 gnd vdd FILL
XNOR2X1_11 Y[17] Y[16] gnd AND2X2_5/A vdd NOR2X1
XINVX1_14 INVX1_14/A gnd INVX1_14/Y vdd INVX1
XFILL_6_2 gnd vdd FILL
XFILL_1_0_1 gnd vdd FILL
XNOR2X1_12 Y[18] Y[19] gnd AND2X2_5/B vdd NOR2X1
XFILL_6_3 gnd vdd FILL
XOAI21X1_10 Y[6] OAI21X1_10/B BUFX2_6/Y gnd XOR2X1_4/A vdd OAI21X1
XFILL_1_0_2 gnd vdd FILL
XNOR2X1_13 Y[21] Y[22] gnd INVX1_4/A vdd NOR2X1
XOAI21X1_11 NOR2X1_5/A NOR2X1_5/B BUFX2_7/Y gnd XNOR2X1_5/A vdd OAI21X1
XFILL_4_0_0 gnd vdd FILL
XFILL_4_1 gnd vdd FILL
XNOR2X1_14 Y[20] Y[23] gnd AND2X2_6/B vdd NOR2X1
XOAI21X1_12 INVX1_1/Y INVX1_11/Y XNOR2X1_5/A gnd XNOR2X1_6/A vdd OAI21X1
XFILL_4_0_1 gnd vdd FILL
XNOR2X1_15 NOR2X1_15/A NOR2X1_15/B gnd NOR2X1_15/Y vdd NOR2X1
XFILL_4_0_2 gnd vdd FILL
XOAI21X1_13 Y[10] OAI21X1_13/B INVX1_1/A gnd XOR2X1_6/A vdd OAI21X1
XNOR2X1_16 Y[24] Y[25] gnd INVX1_2/A vdd NOR2X1
XFILL_2_1_0 gnd vdd FILL
XOAI21X1_14 NOR2X1_10/A NOR3X1_2/A BUFX2_6/Y gnd XOR2X1_7/A vdd OAI21X1
XINVX1_1 INVX1_1/A gnd INVX1_1/Y vdd INVX1
XXNOR2X1_1 XNOR2X1_1/A Y[16] gnd XNOR2X1_1/Y vdd XNOR2X1
XNOR2X1_17 OR2X2_1/Y OR2X2_2/B gnd INVX1_3/A vdd NOR2X1
XAND2X2_1 NOR2X1_1/Y NOR2X1_2/Y gnd AND2X2_1/Y vdd AND2X2
XFILL_2_1 gnd vdd FILL
XFILL_2_1_1 gnd vdd FILL
XOAI21X1_15 Y[12] OAI21X1_16/B BUFX2_7/Y gnd XOR2X1_8/A vdd OAI21X1
XINVX1_2 INVX1_2/A gnd OR2X2_2/B vdd INVX1
XXNOR2X1_2 XNOR2X1_2/A Y[19] gnd XNOR2X1_2/Y vdd XNOR2X1
XAND2X2_2 NOR2X1_3/Y NOR2X1_4/Y gnd AND2X2_2/Y vdd AND2X2
XNOR2X1_18 Y[30] Y[29] gnd AND2X2_9/A vdd NOR2X1
XFILL_2_2 gnd vdd FILL
XFILL_2_1_2 gnd vdd FILL
XOAI21X1_16 INVX1_13/Y OAI21X1_16/B BUFX2_8/Y gnd XNOR2X1_7/A vdd OAI21X1
XOR2X2_1 Y[26] Y[27] gnd OR2X2_1/Y vdd OR2X2
XXNOR2X1_3 OR2X2_2/A Y[24] gnd XNOR2X1_3/Y vdd XNOR2X1
XINVX1_3 INVX1_3/A gnd INVX1_3/Y vdd INVX1
XFILL_5_1_0 gnd vdd FILL
XNOR2X1_19 NOR3X1_2/A NOR3X1_2/B gnd NOR2X1_19/Y vdd NOR2X1
XFILL_2_3 gnd vdd FILL
XAND2X2_3 NOR2X1_6/Y NOR2X1_7/Y gnd AND2X2_3/Y vdd AND2X2
XOAI22X1_1 NOR3X1_3/Y OAI22X1_1/B NOR3X1_1/Y OAI22X1_1/D gnd OAI22X1_1/Y vdd OAI22X1
XOAI21X1_17 INVX1_1/Y INVX1_12/Y XNOR2X1_7/A gnd XNOR2X1_8/A vdd OAI21X1
XOR2X2_2 OR2X2_2/A OR2X2_2/B gnd OR2X2_2/Y vdd OR2X2
XFILL_5_1_1 gnd vdd FILL
XINVX1_4 INVX1_4/A gnd INVX1_4/Y vdd INVX1
XXNOR2X1_4 XNOR2X1_4/A Y[20] gnd XNOR2X1_4/Y vdd XNOR2X1
XAND2X2_4 NOR2X1_8/Y NOR2X1_9/Y gnd AND2X2_4/Y vdd AND2X2
XNAND2X1_20 AND2X2_3/Y NOR2X1_5/Y gnd OAI21X1_16/B vdd NAND2X1
XXNOR2X1_5 XNOR2X1_5/A INVX1_11/Y gnd NOR3X1_8/B vdd XNOR2X1
XINVX1_5 Y[20] gnd INVX1_5/Y vdd INVX1
XOR2X2_3 OR2X2_3/A OR2X2_3/B gnd OR2X2_3/Y vdd OR2X2
.ends

