magic
tech scmos
magscale 1 2
timestamp 1646624542
<< checkpaint >>
rect -76 -66 124 270
<< nwell >>
rect -16 96 64 210
<< ntransistor >>
rect 14 12 18 52
rect 24 12 28 52
<< ptransistor >>
rect 14 148 18 188
rect 30 148 34 188
<< ndiffusion >>
rect 4 51 14 52
rect 12 13 14 51
rect 4 12 14 13
rect 18 12 24 52
rect 28 51 38 52
rect 28 13 30 51
rect 28 12 38 13
<< pdiffusion >>
rect 4 187 14 188
rect 12 149 14 187
rect 4 148 14 149
rect 18 187 30 188
rect 18 149 20 187
rect 28 149 30 187
rect 18 148 30 149
rect 34 187 44 188
rect 34 149 36 187
rect 34 148 44 149
<< ndcontact >>
rect 4 13 12 51
rect 30 13 38 51
<< pdcontact >>
rect 4 149 12 187
rect 20 149 28 187
rect 36 149 44 187
<< psubstratepcontact >>
rect -4 -4 4 4
rect 28 -4 36 4
<< nsubstratencontact >>
rect -4 196 4 204
rect 28 196 36 204
<< polysilicon >>
rect 14 188 18 192
rect 30 188 34 192
rect 14 66 18 148
rect 12 58 18 66
rect 30 122 34 148
rect 30 114 36 122
rect 30 58 34 114
rect 14 52 18 58
rect 24 54 34 58
rect 24 52 28 54
rect 14 8 18 12
rect 24 8 28 12
<< polycontact >>
rect 4 58 12 66
rect 36 114 44 122
<< metal1 >>
rect -4 204 52 206
rect 4 196 28 204
rect 36 196 52 204
rect -4 194 52 196
rect 4 187 12 194
rect 4 148 12 149
rect 20 187 28 188
rect 4 66 12 74
rect 20 52 28 149
rect 36 187 44 194
rect 36 148 44 149
rect 36 106 44 114
rect 4 51 12 52
rect 20 51 38 52
rect 20 46 30 51
rect 4 6 12 13
rect 30 12 38 13
rect -4 4 52 6
rect 4 -4 28 4
rect 36 -4 52 4
rect -4 -6 52 -4
<< m1p >>
rect 36 106 44 114
rect 20 86 28 94
rect 4 66 12 74
<< labels >>
rlabel metal1 8 200 8 200 4 vdd
rlabel metal1 24 90 24 90 4 Y
rlabel metal1 8 0 8 0 4 gnd
rlabel metal1 8 70 8 70 4 A
rlabel metal1 40 110 40 110 4 B
<< end >>
