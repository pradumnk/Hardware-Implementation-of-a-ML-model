magic
tech scmos
magscale 1 2
timestamp 1651685240
<< metal1 >>
rect 1240 1406 1246 1414
rect 1254 1406 1260 1414
rect 1268 1406 1274 1414
rect 1282 1406 1288 1414
rect 445 1357 467 1363
rect 660 1357 691 1363
rect 701 1357 723 1363
rect 909 1357 931 1363
rect 269 1337 323 1343
rect 477 1337 572 1343
rect 893 1337 908 1343
rect 132 1317 147 1323
rect 157 1317 172 1323
rect 317 1317 332 1323
rect 1016 1316 1020 1324
rect 1053 1323 1059 1336
rect 1053 1317 1075 1323
rect 1085 1317 1100 1323
rect 1284 1317 1331 1323
rect 356 1236 358 1244
rect 488 1206 494 1214
rect 502 1206 508 1214
rect 516 1206 522 1214
rect 530 1206 536 1214
rect 964 1176 966 1184
rect 52 1097 67 1103
rect 612 1097 643 1103
rect 804 1097 819 1103
rect 989 1103 995 1123
rect 1460 1114 1464 1122
rect 989 1097 1011 1103
rect 1069 1097 1132 1103
rect 1005 1084 1011 1097
rect 1181 1097 1212 1103
rect 1741 1097 1788 1103
rect 365 1077 380 1083
rect 852 1077 867 1083
rect 877 1077 892 1083
rect 932 1077 947 1083
rect 1101 1077 1116 1083
rect 1716 1077 1731 1083
rect 420 1056 428 1064
rect 893 1057 899 1076
rect 1188 1057 1203 1063
rect 1213 1057 1244 1063
rect 1364 1057 1379 1063
rect 1492 1057 1507 1063
rect 328 1036 332 1044
rect 1240 1006 1246 1014
rect 1254 1006 1260 1014
rect 1268 1006 1274 1014
rect 1282 1006 1288 1014
rect 724 977 766 983
rect 1028 977 1059 983
rect 1368 976 1372 984
rect 1668 976 1672 984
rect 1773 977 1788 983
rect 813 957 828 963
rect 909 957 947 963
rect 397 943 403 956
rect 381 937 403 943
rect 468 936 472 944
rect 797 937 851 943
rect 868 937 899 943
rect 916 937 963 943
rect 1101 937 1116 943
rect 1229 937 1315 943
rect 1492 937 1507 943
rect 1517 937 1532 943
rect 109 917 147 923
rect 253 917 284 923
rect 344 896 348 904
rect 413 897 435 903
rect 644 897 659 903
rect 1565 897 1580 903
rect 488 806 494 814
rect 502 806 508 814
rect 516 806 522 814
rect 530 806 536 814
rect 74 736 76 744
rect 1261 737 1308 743
rect 468 717 515 723
rect 100 697 115 703
rect 445 697 531 703
rect 445 677 451 697
rect 749 697 787 703
rect 1165 697 1180 703
rect 1684 697 1699 703
rect 712 677 732 683
rect 1053 677 1075 683
rect 116 657 131 663
rect 408 636 412 644
rect 996 636 1000 644
rect 1544 636 1548 644
rect 1240 606 1246 614
rect 1254 606 1260 614
rect 1268 606 1274 614
rect 1282 606 1288 614
rect 122 576 124 584
rect 842 576 844 584
rect 340 557 355 563
rect 717 557 732 563
rect 1549 557 1564 563
rect 141 537 156 543
rect 957 537 988 543
rect 1037 524 1043 543
rect 1373 537 1388 543
rect 1725 537 1740 543
rect 573 517 611 523
rect 621 517 652 523
rect 941 517 972 523
rect 1044 517 1059 523
rect 1252 517 1315 523
rect 1773 517 1788 523
rect 461 497 531 503
rect 260 436 264 444
rect 1444 436 1448 444
rect 1764 436 1766 444
rect 488 406 494 414
rect 502 406 508 414
rect 516 406 522 414
rect 530 406 536 414
rect 228 376 230 384
rect 1204 376 1206 384
rect 772 316 780 324
rect 733 297 764 303
rect 1076 297 1091 303
rect 1213 297 1276 303
rect 1517 297 1619 303
rect 189 277 204 283
rect 189 257 195 277
rect 525 277 604 283
rect 669 277 700 283
rect 989 277 1011 283
rect 1252 277 1283 283
rect 1325 277 1356 283
rect 1421 277 1436 283
rect 1613 277 1619 297
rect 1741 277 1788 283
rect 285 257 312 263
rect 1412 257 1427 263
rect 52 236 62 244
rect 468 236 472 244
rect 580 237 638 243
rect 872 236 876 244
rect 1156 236 1158 244
rect 1650 237 1692 243
rect 1240 206 1246 214
rect 1254 206 1260 214
rect 1268 206 1274 214
rect 1282 206 1288 214
rect 1064 176 1068 184
rect 253 157 268 163
rect 429 157 444 163
rect 877 157 892 163
rect 228 137 259 143
rect 861 137 876 143
rect 93 117 115 123
rect 205 117 252 123
rect 381 117 412 123
rect 1005 123 1011 143
rect 1581 137 1596 143
rect 868 117 915 123
rect 989 117 1036 123
rect 1165 117 1292 123
rect 1565 117 1612 123
rect 488 6 494 14
rect 502 6 508 14
rect 516 6 522 14
rect 530 6 536 14
<< m2contact >>
rect 1246 1406 1254 1414
rect 1260 1406 1268 1414
rect 1274 1406 1282 1414
rect 1356 1376 1364 1384
rect 1404 1376 1412 1384
rect 1452 1376 1460 1384
rect 1500 1376 1508 1384
rect 1548 1376 1556 1384
rect 1596 1376 1604 1384
rect 1644 1376 1652 1384
rect 1692 1376 1700 1384
rect 1740 1376 1748 1384
rect 28 1358 36 1366
rect 204 1356 212 1364
rect 220 1356 228 1364
rect 284 1356 292 1364
rect 300 1356 308 1364
rect 396 1356 404 1364
rect 636 1356 644 1364
rect 652 1356 660 1364
rect 940 1356 948 1364
rect 1100 1356 1108 1364
rect 1132 1356 1140 1364
rect 1244 1356 1252 1364
rect 1436 1358 1444 1366
rect 1532 1358 1540 1366
rect 1580 1358 1588 1366
rect 1628 1358 1636 1366
rect 1676 1358 1684 1366
rect 1724 1358 1732 1366
rect 1788 1356 1796 1364
rect 108 1336 116 1344
rect 172 1336 180 1344
rect 332 1336 340 1344
rect 412 1336 420 1344
rect 572 1336 580 1344
rect 604 1336 612 1344
rect 636 1336 644 1344
rect 748 1336 756 1344
rect 780 1336 788 1344
rect 844 1336 852 1344
rect 876 1336 884 1344
rect 908 1336 916 1344
rect 956 1336 964 1344
rect 1052 1336 1060 1344
rect 1196 1336 1204 1344
rect 1228 1336 1236 1344
rect 44 1316 52 1324
rect 92 1316 100 1324
rect 124 1316 132 1324
rect 172 1316 180 1324
rect 188 1316 196 1324
rect 332 1316 340 1324
rect 348 1316 356 1324
rect 492 1316 500 1324
rect 620 1316 628 1324
rect 732 1316 740 1324
rect 764 1316 772 1324
rect 796 1316 804 1324
rect 828 1316 836 1324
rect 860 1316 868 1324
rect 1020 1316 1028 1324
rect 1100 1316 1108 1324
rect 1212 1316 1220 1324
rect 1276 1316 1284 1324
rect 1372 1316 1380 1324
rect 1420 1316 1428 1324
rect 1468 1316 1476 1324
rect 1516 1316 1524 1324
rect 1564 1316 1572 1324
rect 1612 1316 1620 1324
rect 1660 1316 1668 1324
rect 1708 1316 1716 1324
rect 1756 1316 1764 1324
rect 124 1296 132 1304
rect 236 1296 244 1304
rect 380 1296 388 1304
rect 12 1276 20 1284
rect 60 1236 68 1244
rect 348 1236 356 1244
rect 812 1236 820 1244
rect 1116 1236 1124 1244
rect 1756 1236 1764 1244
rect 494 1206 502 1214
rect 508 1206 516 1214
rect 522 1206 530 1214
rect 956 1176 964 1184
rect 1132 1176 1140 1184
rect 1308 1176 1316 1184
rect 1692 1156 1700 1164
rect 60 1136 68 1144
rect 44 1116 52 1124
rect 140 1116 148 1124
rect 604 1116 612 1124
rect 620 1116 628 1124
rect 684 1116 692 1124
rect 700 1116 708 1124
rect 844 1116 852 1124
rect 44 1096 52 1104
rect 172 1096 180 1104
rect 220 1096 228 1104
rect 380 1096 388 1104
rect 444 1096 452 1104
rect 508 1096 516 1104
rect 604 1096 612 1104
rect 652 1096 660 1104
rect 764 1096 772 1104
rect 796 1096 804 1104
rect 828 1096 836 1104
rect 924 1096 932 1104
rect 956 1096 964 1104
rect 1452 1114 1460 1122
rect 1548 1116 1556 1124
rect 1132 1096 1140 1104
rect 1212 1096 1220 1104
rect 1356 1096 1364 1104
rect 1484 1096 1492 1104
rect 1628 1096 1636 1104
rect 1660 1096 1668 1104
rect 1788 1096 1796 1104
rect 12 1076 20 1084
rect 124 1076 132 1084
rect 156 1076 164 1084
rect 188 1076 196 1084
rect 204 1076 212 1084
rect 268 1076 276 1084
rect 380 1076 388 1084
rect 396 1076 404 1084
rect 428 1076 436 1084
rect 524 1076 532 1084
rect 572 1076 580 1084
rect 588 1076 596 1084
rect 668 1076 676 1084
rect 716 1076 724 1084
rect 780 1076 788 1084
rect 844 1076 852 1084
rect 892 1076 900 1084
rect 924 1076 932 1084
rect 1004 1076 1012 1084
rect 1116 1076 1124 1084
rect 1196 1076 1204 1084
rect 1372 1076 1380 1084
rect 1500 1076 1508 1084
rect 1580 1076 1588 1084
rect 1644 1076 1652 1084
rect 1708 1076 1716 1084
rect 92 1056 100 1064
rect 108 1056 116 1064
rect 428 1056 436 1064
rect 556 1056 564 1064
rect 796 1056 804 1064
rect 908 1056 916 1064
rect 1180 1056 1188 1064
rect 1244 1056 1252 1064
rect 1356 1056 1364 1064
rect 1484 1056 1492 1064
rect 1708 1056 1716 1064
rect 44 1036 52 1044
rect 252 1036 260 1044
rect 332 1036 340 1044
rect 540 1036 548 1044
rect 732 1036 740 1044
rect 1548 1036 1556 1044
rect 1596 1036 1604 1044
rect 1740 1016 1748 1024
rect 1246 1006 1254 1014
rect 1260 1006 1268 1014
rect 1274 1006 1282 1014
rect 28 976 36 984
rect 716 976 724 984
rect 956 976 964 984
rect 1020 976 1028 984
rect 1196 976 1204 984
rect 1372 976 1380 984
rect 1660 976 1668 984
rect 1788 976 1796 984
rect 12 956 20 964
rect 396 956 404 964
rect 828 956 836 964
rect 860 956 868 964
rect 956 956 964 964
rect 1116 956 1124 964
rect 60 936 68 944
rect 220 936 228 944
rect 284 936 292 944
rect 460 936 468 944
rect 604 936 612 944
rect 860 936 868 944
rect 908 936 916 944
rect 1116 936 1124 944
rect 1212 936 1220 944
rect 1404 936 1412 944
rect 1436 936 1444 944
rect 1468 936 1476 944
rect 1484 936 1492 944
rect 1532 936 1540 944
rect 1580 936 1588 944
rect 1628 936 1636 944
rect 1724 936 1732 944
rect 44 916 52 924
rect 76 916 84 924
rect 188 916 196 924
rect 204 916 212 924
rect 236 916 244 924
rect 284 916 292 924
rect 444 916 452 924
rect 556 916 564 924
rect 668 916 676 924
rect 780 916 788 924
rect 876 916 884 924
rect 972 916 980 924
rect 1084 916 1092 924
rect 1148 916 1156 924
rect 1164 916 1172 924
rect 1452 916 1460 924
rect 1740 916 1748 924
rect 156 896 164 904
rect 268 896 276 904
rect 348 896 356 904
rect 588 896 596 904
rect 620 896 628 904
rect 636 896 644 904
rect 1052 896 1060 904
rect 1244 896 1252 904
rect 1420 896 1428 904
rect 1484 896 1492 904
rect 1580 896 1588 904
rect 1612 896 1620 904
rect 460 876 468 884
rect 556 876 564 884
rect 684 876 692 884
rect 572 836 580 844
rect 668 836 676 844
rect 1148 836 1156 844
rect 1548 836 1556 844
rect 1596 836 1604 844
rect 494 806 502 814
rect 508 806 516 814
rect 522 806 530 814
rect 188 776 196 784
rect 236 776 244 784
rect 924 776 932 784
rect 1132 776 1140 784
rect 1212 776 1220 784
rect 1628 776 1636 784
rect 1644 776 1652 784
rect 1724 776 1732 784
rect 1772 776 1780 784
rect 316 756 324 764
rect 828 756 836 764
rect 12 736 20 744
rect 76 736 84 744
rect 172 736 180 744
rect 252 736 260 744
rect 300 736 308 744
rect 700 736 708 744
rect 892 736 900 744
rect 1308 736 1316 744
rect 204 716 212 724
rect 220 716 228 724
rect 332 716 340 724
rect 460 716 468 724
rect 668 716 676 724
rect 732 716 740 724
rect 860 716 868 724
rect 1068 716 1076 724
rect 1404 716 1412 724
rect 1420 716 1428 724
rect 44 696 52 704
rect 60 696 68 704
rect 92 696 100 704
rect 188 696 196 704
rect 236 696 244 704
rect 316 696 324 704
rect 348 676 356 684
rect 540 696 548 704
rect 588 696 596 704
rect 620 696 628 704
rect 652 696 660 704
rect 684 696 692 704
rect 844 696 852 704
rect 876 696 884 704
rect 1100 696 1108 704
rect 1180 696 1188 704
rect 1228 696 1236 704
rect 1356 696 1364 704
rect 1452 696 1460 704
rect 1628 696 1636 704
rect 1676 696 1684 704
rect 1740 696 1748 704
rect 556 676 564 684
rect 604 676 612 684
rect 732 676 740 684
rect 764 676 772 684
rect 796 676 804 684
rect 828 676 836 684
rect 956 676 964 684
rect 1116 676 1124 684
rect 1324 676 1332 684
rect 1372 676 1380 684
rect 1436 676 1444 684
rect 1468 676 1476 684
rect 1484 676 1492 684
rect 1580 676 1588 684
rect 28 654 36 662
rect 92 656 100 664
rect 108 656 116 664
rect 140 656 148 664
rect 572 656 580 664
rect 636 656 644 664
rect 940 656 948 664
rect 1596 656 1604 664
rect 1660 654 1668 662
rect 412 636 420 644
rect 732 636 740 644
rect 892 636 900 644
rect 924 636 932 644
rect 988 636 996 644
rect 1132 636 1140 644
rect 1212 636 1220 644
rect 1404 636 1412 644
rect 1548 636 1556 644
rect 1612 636 1620 644
rect 92 616 100 624
rect 1246 606 1254 614
rect 1260 606 1268 614
rect 1274 606 1282 614
rect 1740 596 1748 604
rect 124 576 132 584
rect 204 576 212 584
rect 684 576 692 584
rect 844 576 852 584
rect 956 576 964 584
rect 1116 576 1124 584
rect 1756 576 1764 584
rect 28 558 36 566
rect 332 556 340 564
rect 364 556 372 564
rect 380 556 388 564
rect 444 556 452 564
rect 732 556 740 564
rect 764 556 772 564
rect 972 556 980 564
rect 1388 556 1396 564
rect 1564 556 1572 564
rect 1740 556 1748 564
rect 60 536 68 544
rect 156 536 164 544
rect 220 536 228 544
rect 316 536 324 544
rect 412 536 420 544
rect 588 536 596 544
rect 652 536 660 544
rect 860 536 868 544
rect 988 536 996 544
rect 1100 536 1108 544
rect 1148 536 1156 544
rect 1196 536 1204 544
rect 1340 536 1348 544
rect 1388 536 1396 544
rect 1404 536 1412 544
rect 1500 536 1508 544
rect 1548 536 1556 544
rect 1740 536 1748 544
rect 44 516 52 524
rect 92 516 100 524
rect 172 516 180 524
rect 332 516 340 524
rect 396 516 404 524
rect 428 516 436 524
rect 540 516 548 524
rect 652 516 660 524
rect 732 516 740 524
rect 748 516 756 524
rect 812 516 820 524
rect 972 516 980 524
rect 1036 516 1044 524
rect 1084 516 1092 524
rect 1244 516 1252 524
rect 1356 516 1364 524
rect 1564 516 1572 524
rect 1644 516 1652 524
rect 1692 516 1700 524
rect 1788 516 1796 524
rect 108 496 116 504
rect 636 496 644 504
rect 684 496 692 504
rect 828 496 836 504
rect 1004 496 1012 504
rect 1116 496 1124 504
rect 1164 496 1172 504
rect 1612 496 1620 504
rect 12 476 20 484
rect 556 476 564 484
rect 1212 476 1220 484
rect 1676 476 1684 484
rect 540 456 548 464
rect 252 436 260 444
rect 700 436 708 444
rect 780 436 788 444
rect 1020 436 1028 444
rect 1180 436 1188 444
rect 1436 436 1444 444
rect 1756 436 1764 444
rect 494 406 502 414
rect 508 406 516 414
rect 522 406 530 414
rect 220 376 228 384
rect 1196 376 1204 384
rect 316 336 324 344
rect 252 316 260 324
rect 348 316 356 324
rect 764 316 772 324
rect 796 316 804 324
rect 1052 316 1060 324
rect 1116 316 1124 324
rect 1164 316 1172 324
rect 1324 316 1332 324
rect 76 296 84 304
rect 220 296 228 304
rect 332 296 340 304
rect 412 296 420 304
rect 652 296 660 304
rect 764 296 772 304
rect 956 296 964 304
rect 1020 296 1028 304
rect 1036 296 1044 304
rect 1068 296 1076 304
rect 1276 296 1284 304
rect 1292 296 1300 304
rect 1404 296 1412 304
rect 92 276 100 284
rect 172 276 180 284
rect 108 256 116 264
rect 204 276 212 284
rect 380 276 388 284
rect 396 276 404 284
rect 428 276 436 284
rect 604 276 612 284
rect 700 276 708 284
rect 748 276 756 284
rect 812 276 820 284
rect 908 276 916 284
rect 1068 276 1076 284
rect 1100 276 1108 284
rect 1132 276 1140 284
rect 1244 276 1252 284
rect 1356 276 1364 284
rect 1436 276 1444 284
rect 1468 276 1476 284
rect 1564 276 1572 284
rect 1628 296 1636 304
rect 1708 296 1716 304
rect 1788 276 1796 284
rect 268 256 276 264
rect 364 256 372 264
rect 684 256 692 264
rect 716 256 724 264
rect 972 256 980 264
rect 1180 256 1188 264
rect 1404 256 1412 264
rect 1596 256 1604 264
rect 1724 254 1732 262
rect 44 236 52 244
rect 140 236 148 244
rect 460 236 468 244
rect 572 236 580 244
rect 876 236 884 244
rect 924 236 932 244
rect 1148 236 1156 244
rect 1420 236 1428 244
rect 1692 236 1700 244
rect 1246 206 1254 214
rect 1260 206 1268 214
rect 1274 206 1282 214
rect 252 176 260 184
rect 428 176 436 184
rect 668 176 676 184
rect 732 176 740 184
rect 860 176 868 184
rect 972 176 980 184
rect 1068 176 1076 184
rect 1676 176 1684 184
rect 268 156 276 164
rect 444 156 452 164
rect 652 156 660 164
rect 892 156 900 164
rect 956 156 964 164
rect 1356 156 1364 164
rect 1580 156 1588 164
rect 60 136 68 144
rect 156 136 164 144
rect 220 136 228 144
rect 428 136 436 144
rect 716 136 724 144
rect 764 136 772 144
rect 876 136 884 144
rect 44 116 52 124
rect 140 116 148 124
rect 252 116 260 124
rect 268 116 276 124
rect 412 116 420 124
rect 444 116 452 124
rect 572 116 580 124
rect 620 116 628 124
rect 636 116 644 124
rect 700 116 708 124
rect 844 116 852 124
rect 860 116 868 124
rect 1100 136 1108 144
rect 1116 136 1124 144
rect 1212 136 1220 144
rect 1324 136 1332 144
rect 1356 136 1364 144
rect 1548 136 1556 144
rect 1596 136 1604 144
rect 1724 136 1732 144
rect 1036 116 1044 124
rect 1292 116 1300 124
rect 1340 116 1348 124
rect 1404 116 1412 124
rect 1452 116 1460 124
rect 1612 116 1620 124
rect 1628 116 1636 124
rect 1708 116 1716 124
rect 1772 116 1780 124
rect 732 96 740 104
rect 12 76 20 84
rect 172 36 180 44
rect 348 36 356 44
rect 604 36 612 44
rect 940 36 948 44
rect 1436 36 1444 44
rect 1484 36 1492 44
rect 1660 36 1668 44
rect 1740 36 1748 44
rect 494 6 502 14
rect 508 6 516 14
rect 522 6 530 14
<< metal2 >>
rect 36 1358 51 1363
rect 29 1357 51 1358
rect 45 1324 51 1357
rect 13 1284 19 1296
rect 109 1284 115 1336
rect 189 1324 195 1443
rect 221 1437 243 1443
rect 221 1364 227 1437
rect 221 1344 227 1356
rect 189 1304 195 1316
rect 61 1163 67 1236
rect 61 1157 83 1163
rect 61 1124 67 1136
rect 52 1117 60 1123
rect 20 1077 35 1083
rect 29 1064 35 1077
rect 29 984 35 1056
rect 45 964 51 1036
rect 13 944 19 956
rect 77 944 83 1157
rect 141 1104 147 1116
rect 221 1104 227 1116
rect 157 1064 163 1076
rect 93 1044 99 1056
rect 93 964 99 1036
rect 173 924 179 1096
rect 269 1084 275 1336
rect 285 1324 291 1356
rect 397 1344 403 1356
rect 413 1344 419 1443
rect 637 1364 643 1443
rect 861 1404 867 1443
rect 285 1284 291 1316
rect 349 1304 355 1316
rect 413 1304 419 1336
rect 493 1324 499 1356
rect 621 1343 627 1356
rect 653 1344 659 1356
rect 749 1344 755 1376
rect 621 1337 636 1343
rect 349 1144 355 1236
rect 381 1104 387 1276
rect 488 1206 494 1214
rect 502 1206 508 1214
rect 516 1206 522 1214
rect 530 1206 536 1214
rect 381 1084 387 1096
rect 429 1084 435 1136
rect 445 1084 451 1096
rect 205 1044 211 1076
rect 189 924 195 1036
rect 253 1024 259 1036
rect 333 984 339 1036
rect 45 904 51 916
rect 77 904 83 916
rect 237 904 243 916
rect 253 883 259 936
rect 237 877 259 883
rect 189 784 195 876
rect 61 704 67 716
rect 189 704 195 736
rect 221 724 227 816
rect 237 784 243 877
rect 45 663 51 696
rect 29 662 51 663
rect 36 657 51 662
rect 93 644 99 656
rect 36 558 51 563
rect 29 557 51 558
rect 45 524 51 557
rect 93 524 99 616
rect 109 524 115 656
rect 125 584 131 636
rect 205 624 211 716
rect 221 603 227 716
rect 237 624 243 696
rect 269 684 275 896
rect 285 844 291 916
rect 381 884 387 1076
rect 397 1064 403 1076
rect 509 1064 515 1096
rect 525 1084 531 1096
rect 573 1084 579 1336
rect 605 1324 611 1336
rect 829 1324 835 1336
rect 621 1284 627 1316
rect 733 1304 739 1316
rect 797 1304 803 1316
rect 845 1284 851 1336
rect 605 1124 611 1136
rect 685 1124 691 1276
rect 653 1084 659 1096
rect 685 1083 691 1116
rect 676 1077 691 1083
rect 541 1004 547 1036
rect 557 984 563 1056
rect 461 924 467 936
rect 445 824 451 916
rect 477 883 483 936
rect 468 877 483 883
rect 541 883 547 976
rect 557 904 563 916
rect 573 884 579 1076
rect 669 1024 675 1076
rect 717 1064 723 1076
rect 781 1064 787 1076
rect 541 877 556 883
rect 445 784 451 816
rect 488 806 494 814
rect 502 806 508 814
rect 516 806 522 814
rect 530 806 536 814
rect 573 804 579 836
rect 205 597 227 603
rect 205 584 211 597
rect 301 584 307 736
rect 317 724 323 756
rect 589 744 595 896
rect 605 784 611 936
rect 637 904 643 1016
rect 717 984 723 1016
rect 685 884 691 956
rect 733 924 739 1036
rect 781 864 787 916
rect 317 624 323 696
rect 157 544 163 556
rect 221 544 227 576
rect 333 564 339 716
rect 349 684 355 696
rect 317 524 323 536
rect 333 524 339 536
rect 109 504 115 516
rect 333 504 339 516
rect 13 484 19 496
rect 221 384 227 476
rect 253 324 259 436
rect 317 344 323 356
rect 349 324 355 336
rect 93 284 99 316
rect 365 304 371 556
rect 381 384 387 556
rect 413 544 419 616
rect 429 524 435 576
rect 445 504 451 556
rect 413 364 419 456
rect 413 304 419 356
rect 461 344 467 716
rect 541 704 547 716
rect 605 684 611 756
rect 621 704 627 796
rect 637 704 643 776
rect 669 764 675 836
rect 669 724 675 736
rect 701 724 707 736
rect 797 724 803 1056
rect 717 717 732 723
rect 717 684 723 717
rect 813 683 819 1236
rect 829 1104 835 1196
rect 861 1144 867 1316
rect 845 1104 851 1116
rect 829 964 835 1096
rect 861 1084 867 1136
rect 877 963 883 1336
rect 893 1084 899 1443
rect 925 1363 931 1443
rect 925 1357 940 1363
rect 925 1204 931 1357
rect 1053 1344 1059 1443
rect 1101 1437 1123 1443
rect 1101 1364 1107 1437
rect 1240 1406 1246 1414
rect 1254 1406 1260 1414
rect 1268 1406 1274 1414
rect 1282 1406 1288 1414
rect 1325 1404 1331 1443
rect 1373 1404 1379 1443
rect 1421 1404 1427 1443
rect 1485 1437 1507 1443
rect 1533 1437 1555 1443
rect 1581 1437 1603 1443
rect 1629 1437 1651 1443
rect 1677 1437 1699 1443
rect 1725 1437 1747 1443
rect 1357 1384 1363 1396
rect 1405 1384 1411 1396
rect 1453 1384 1459 1396
rect 1501 1384 1507 1437
rect 1549 1384 1555 1437
rect 1597 1384 1603 1437
rect 1645 1384 1651 1437
rect 1693 1384 1699 1437
rect 1741 1384 1747 1437
rect 1757 1437 1779 1443
rect 1789 1437 1811 1443
rect 1421 1358 1436 1363
rect 1517 1358 1532 1363
rect 1565 1358 1580 1363
rect 1613 1358 1628 1363
rect 1661 1358 1676 1363
rect 1709 1358 1724 1363
rect 1421 1357 1443 1358
rect 1517 1357 1539 1358
rect 1565 1357 1587 1358
rect 1613 1357 1635 1358
rect 1661 1357 1683 1358
rect 1709 1357 1731 1358
rect 957 1184 963 1336
rect 1197 1324 1203 1336
rect 925 984 931 1076
rect 957 984 963 1076
rect 1005 1043 1011 1076
rect 1005 1037 1027 1043
rect 1021 984 1027 1037
rect 868 957 883 963
rect 909 924 915 936
rect 845 704 851 736
rect 861 724 867 836
rect 877 704 883 776
rect 893 744 899 756
rect 909 684 915 916
rect 925 784 931 976
rect 957 804 963 956
rect 1085 924 1091 936
rect 973 904 979 916
rect 1101 824 1107 1316
rect 1117 1104 1123 1236
rect 1133 1184 1139 1296
rect 1213 1104 1219 1316
rect 1117 1084 1123 1096
rect 1133 1084 1139 1096
rect 1213 1063 1219 1096
rect 1245 1064 1251 1356
rect 1421 1324 1427 1357
rect 1517 1324 1523 1357
rect 1565 1324 1571 1357
rect 1613 1324 1619 1357
rect 1661 1324 1667 1357
rect 1709 1324 1715 1357
rect 1757 1324 1763 1437
rect 1789 1364 1795 1437
rect 1309 1184 1315 1316
rect 1373 1304 1379 1316
rect 1549 1104 1555 1116
rect 1661 1104 1667 1116
rect 1757 1104 1763 1236
rect 1789 1104 1795 1116
rect 1197 1057 1219 1063
rect 1181 1004 1187 1056
rect 1197 984 1203 1057
rect 1240 1006 1246 1014
rect 1254 1006 1260 1014
rect 1268 1006 1274 1014
rect 1282 1006 1288 1014
rect 1373 984 1379 1076
rect 1501 1064 1507 1076
rect 1117 944 1123 956
rect 1437 944 1443 956
rect 1117 924 1123 936
rect 1149 924 1155 936
rect 1069 724 1075 736
rect 813 677 828 683
rect 557 664 563 676
rect 644 657 659 663
rect 573 644 579 656
rect 589 544 595 556
rect 653 544 659 657
rect 685 584 691 676
rect 733 564 739 636
rect 765 564 771 576
rect 541 524 547 536
rect 557 484 563 516
rect 653 504 659 516
rect 637 444 643 496
rect 488 406 494 414
rect 502 406 508 414
rect 516 406 522 414
rect 530 406 536 414
rect 45 124 51 236
rect 109 184 115 256
rect 141 144 147 236
rect 157 144 163 296
rect 221 284 227 296
rect 205 264 211 276
rect 365 264 371 296
rect 397 284 403 296
rect 429 284 435 316
rect 653 304 659 416
rect 612 277 627 283
rect 157 124 163 136
rect 253 124 259 176
rect 269 164 275 176
rect 13 84 19 96
rect 173 -17 179 36
rect 173 -23 195 -17
rect 349 -23 355 36
rect 365 -17 371 256
rect 429 163 435 176
rect 445 164 451 176
rect 413 157 435 163
rect 413 124 419 157
rect 461 144 467 236
rect 573 124 579 236
rect 621 124 627 277
rect 653 164 659 256
rect 669 184 675 456
rect 701 284 707 436
rect 685 184 691 256
rect 733 184 739 516
rect 797 484 803 676
rect 813 524 819 636
rect 845 584 851 676
rect 941 664 947 716
rect 1101 704 1107 796
rect 1133 784 1139 896
rect 861 524 867 536
rect 829 464 835 496
rect 749 284 755 356
rect 765 284 771 296
rect 605 24 611 36
rect 488 6 494 14
rect 502 6 508 14
rect 516 6 522 14
rect 530 6 536 14
rect 365 -23 387 -17
rect 573 -23 579 16
rect 621 -17 627 116
rect 605 -23 627 -17
rect 653 -23 659 156
rect 717 144 723 156
rect 765 144 771 156
rect 781 144 787 436
rect 925 364 931 636
rect 797 304 803 316
rect 957 304 963 576
rect 973 564 979 596
rect 989 544 995 636
rect 1117 584 1123 676
rect 1133 584 1139 636
rect 1149 563 1155 836
rect 1165 644 1171 916
rect 1213 904 1219 936
rect 1245 904 1251 916
rect 1405 864 1411 936
rect 1421 844 1427 896
rect 1469 864 1475 936
rect 1533 844 1539 936
rect 1549 924 1555 1036
rect 1597 943 1603 1036
rect 1661 984 1667 1056
rect 1629 944 1635 956
rect 1588 937 1603 943
rect 1581 904 1587 936
rect 1741 924 1747 1016
rect 1789 984 1795 1016
rect 1165 584 1171 636
rect 1197 564 1203 816
rect 1213 784 1219 836
rect 1421 724 1427 736
rect 1549 724 1555 836
rect 1597 804 1603 836
rect 1453 704 1459 716
rect 1581 684 1587 736
rect 1380 677 1395 683
rect 1325 664 1331 676
rect 1149 557 1171 563
rect 1101 544 1107 556
rect 1133 543 1139 556
rect 1165 544 1171 557
rect 1197 544 1203 556
rect 1133 537 1148 543
rect 973 484 979 516
rect 1005 504 1011 536
rect 1117 504 1123 516
rect 1165 504 1171 536
rect 1213 504 1219 636
rect 1240 606 1246 614
rect 1254 606 1260 614
rect 1268 606 1274 614
rect 1282 606 1288 614
rect 1245 524 1251 576
rect 973 424 979 476
rect 1021 324 1027 436
rect 1117 384 1123 496
rect 1053 324 1059 336
rect 1021 304 1027 316
rect 1053 304 1059 316
rect 1069 304 1075 316
rect 1133 304 1139 496
rect 1181 323 1187 436
rect 1325 324 1331 656
rect 1389 564 1395 677
rect 1469 664 1475 676
rect 1597 664 1603 776
rect 1613 683 1619 896
rect 1629 784 1635 896
rect 1645 784 1651 876
rect 1789 864 1795 956
rect 1725 784 1731 796
rect 1629 704 1635 736
rect 1613 677 1635 683
rect 1405 544 1411 636
rect 1469 584 1475 656
rect 1501 544 1507 576
rect 1549 544 1555 636
rect 1572 557 1587 563
rect 1341 524 1347 536
rect 1357 484 1363 516
rect 1172 317 1187 323
rect 1181 304 1187 317
rect 909 284 915 296
rect 1133 284 1139 296
rect 861 124 867 176
rect 877 144 883 236
rect 893 164 899 176
rect 733 104 739 116
rect 925 -17 931 236
rect 957 164 963 276
rect 973 184 979 256
rect 973 164 979 176
rect 957 44 963 156
rect 1101 144 1107 276
rect 1181 264 1187 276
rect 1149 184 1155 236
rect 1117 144 1123 176
rect 1213 144 1219 276
rect 1277 264 1283 296
rect 1240 206 1246 214
rect 1254 206 1260 214
rect 1268 206 1274 214
rect 1282 206 1288 214
rect 941 24 947 36
rect 925 -23 947 -17
rect 973 -23 979 16
rect 1005 -23 1011 36
rect 1037 -17 1043 116
rect 1037 -23 1059 -17
rect 1213 -23 1219 136
rect 1293 124 1299 136
rect 1325 124 1331 136
rect 1341 124 1347 476
rect 1405 304 1411 516
rect 1437 284 1443 436
rect 1565 264 1571 276
rect 1405 244 1411 256
rect 1357 164 1363 236
rect 1421 124 1427 236
rect 1549 124 1555 136
rect 1437 24 1443 36
rect 1405 -23 1411 16
rect 1485 -17 1491 36
rect 1565 24 1571 256
rect 1581 244 1587 557
rect 1613 524 1619 636
rect 1629 464 1635 677
rect 1677 663 1683 696
rect 1661 662 1683 663
rect 1668 657 1683 662
rect 1741 604 1747 696
rect 1757 584 1763 836
rect 1773 784 1779 816
rect 1741 564 1747 576
rect 1645 524 1651 536
rect 1789 524 1795 856
rect 1693 504 1699 516
rect 1597 244 1603 256
rect 1581 164 1587 236
rect 1597 144 1603 156
rect 1613 124 1619 296
rect 1677 184 1683 456
rect 1709 263 1715 296
rect 1709 262 1731 263
rect 1709 257 1724 262
rect 1693 224 1699 236
rect 1709 124 1715 236
rect 1757 144 1763 436
rect 1789 284 1795 296
rect 1773 124 1779 216
rect 1469 -23 1491 -17
rect 1517 -23 1523 16
rect 1661 -17 1667 36
rect 1645 -23 1667 -17
rect 1741 -17 1747 36
rect 1741 -23 1763 -17
<< m3contact >>
rect 172 1336 180 1344
rect 92 1316 100 1324
rect 12 1296 20 1304
rect 204 1356 212 1364
rect 300 1356 308 1364
rect 220 1336 228 1344
rect 268 1336 276 1344
rect 124 1316 132 1324
rect 172 1316 180 1324
rect 124 1296 132 1304
rect 188 1296 196 1304
rect 236 1296 244 1304
rect 108 1276 116 1284
rect 60 1116 68 1124
rect 44 1096 52 1104
rect 28 1056 36 1064
rect 44 956 52 964
rect 220 1116 228 1124
rect 140 1096 148 1104
rect 124 1076 132 1084
rect 108 1056 116 1064
rect 156 1056 164 1064
rect 92 1036 100 1044
rect 92 956 100 964
rect 12 936 20 944
rect 60 936 68 944
rect 76 936 84 944
rect 860 1396 868 1404
rect 748 1376 756 1384
rect 492 1356 500 1364
rect 620 1356 628 1364
rect 332 1336 340 1344
rect 396 1336 404 1344
rect 284 1316 292 1324
rect 332 1316 340 1324
rect 652 1336 660 1344
rect 780 1336 788 1344
rect 828 1336 836 1344
rect 492 1316 500 1324
rect 348 1296 356 1304
rect 380 1296 388 1304
rect 412 1296 420 1304
rect 284 1276 292 1284
rect 380 1276 388 1284
rect 348 1136 356 1144
rect 494 1206 502 1214
rect 508 1206 516 1214
rect 522 1206 530 1214
rect 428 1136 436 1144
rect 524 1096 532 1104
rect 188 1076 196 1084
rect 444 1076 452 1084
rect 188 1036 196 1044
rect 204 1036 212 1044
rect 252 1016 260 1024
rect 332 976 340 984
rect 220 936 228 944
rect 252 936 260 944
rect 284 936 292 944
rect 172 916 180 924
rect 204 916 212 924
rect 44 896 52 904
rect 76 896 84 904
rect 156 896 164 904
rect 236 896 244 904
rect 188 876 196 884
rect 220 816 228 824
rect 12 736 20 744
rect 76 736 84 744
rect 172 736 180 744
rect 188 736 196 744
rect 60 716 68 724
rect 252 736 260 744
rect 92 696 100 704
rect 140 656 148 664
rect 92 636 100 644
rect 60 536 68 544
rect 124 636 132 644
rect 204 616 212 624
rect 348 896 356 904
rect 604 1316 612 1324
rect 764 1316 772 1324
rect 732 1296 740 1304
rect 796 1296 804 1304
rect 860 1316 868 1324
rect 620 1276 628 1284
rect 684 1276 692 1284
rect 844 1276 852 1284
rect 604 1136 612 1144
rect 620 1116 628 1124
rect 700 1116 708 1124
rect 604 1096 612 1104
rect 588 1076 596 1084
rect 652 1076 660 1084
rect 764 1096 772 1104
rect 796 1096 804 1104
rect 396 1056 404 1064
rect 428 1056 436 1064
rect 508 1056 516 1064
rect 540 996 548 1004
rect 540 976 548 984
rect 556 976 564 984
rect 396 956 404 964
rect 476 936 484 944
rect 460 916 468 924
rect 380 876 388 884
rect 284 836 292 844
rect 556 896 564 904
rect 716 1056 724 1064
rect 780 1056 788 1064
rect 636 1016 644 1024
rect 668 1016 676 1024
rect 716 1016 724 1024
rect 572 876 580 884
rect 444 816 452 824
rect 494 806 502 814
rect 508 806 516 814
rect 522 806 530 814
rect 572 796 580 804
rect 444 776 452 784
rect 300 736 308 744
rect 268 676 276 684
rect 236 616 244 624
rect 684 956 692 964
rect 668 916 676 924
rect 620 896 628 904
rect 732 916 740 924
rect 684 876 692 884
rect 780 856 788 864
rect 620 796 628 804
rect 604 776 612 784
rect 604 756 612 764
rect 588 736 596 744
rect 316 716 324 724
rect 540 716 548 724
rect 316 616 324 624
rect 220 576 228 584
rect 300 576 308 584
rect 156 556 164 564
rect 348 696 356 704
rect 412 636 420 644
rect 412 616 420 624
rect 332 556 340 564
rect 364 556 372 564
rect 220 536 228 544
rect 332 536 340 544
rect 108 516 116 524
rect 172 516 180 524
rect 316 516 324 524
rect 12 496 20 504
rect 332 496 340 504
rect 220 476 228 484
rect 316 356 324 364
rect 348 336 356 344
rect 92 316 100 324
rect 252 316 260 324
rect 76 296 84 304
rect 428 576 436 584
rect 412 536 420 544
rect 396 516 404 524
rect 428 516 436 524
rect 444 496 452 504
rect 412 456 420 464
rect 380 376 388 384
rect 412 356 420 364
rect 588 696 596 704
rect 636 776 644 784
rect 668 756 676 764
rect 668 736 676 744
rect 700 716 708 724
rect 636 696 644 704
rect 652 696 660 704
rect 684 696 692 704
rect 796 716 804 724
rect 684 676 692 684
rect 716 676 724 684
rect 732 676 740 684
rect 764 676 772 684
rect 828 1196 836 1204
rect 860 1136 868 1144
rect 844 1096 852 1104
rect 844 1076 852 1084
rect 860 1076 868 1084
rect 860 956 868 964
rect 908 1336 916 1344
rect 1246 1406 1254 1414
rect 1260 1406 1268 1414
rect 1274 1406 1282 1414
rect 1324 1396 1332 1404
rect 1356 1396 1364 1404
rect 1372 1396 1380 1404
rect 1404 1396 1412 1404
rect 1420 1396 1428 1404
rect 1452 1396 1460 1404
rect 1100 1356 1108 1364
rect 1132 1356 1140 1364
rect 1228 1336 1236 1344
rect 924 1196 932 1204
rect 1020 1316 1028 1324
rect 1196 1316 1204 1324
rect 924 1096 932 1104
rect 956 1096 964 1104
rect 956 1076 964 1084
rect 908 1056 916 1064
rect 924 976 932 984
rect 860 936 868 944
rect 876 916 884 924
rect 908 916 916 924
rect 860 836 868 844
rect 828 756 836 764
rect 844 736 852 744
rect 876 776 884 784
rect 892 756 900 764
rect 1084 936 1092 944
rect 972 896 980 904
rect 1052 896 1060 904
rect 1132 1296 1140 1304
rect 1116 1096 1124 1104
rect 1212 1096 1220 1104
rect 1132 1076 1140 1084
rect 1196 1076 1204 1084
rect 1276 1316 1284 1324
rect 1308 1316 1316 1324
rect 1468 1316 1476 1324
rect 1372 1296 1380 1304
rect 1692 1156 1700 1164
rect 1452 1122 1460 1124
rect 1452 1116 1460 1122
rect 1660 1116 1668 1124
rect 1788 1116 1796 1124
rect 1356 1096 1364 1104
rect 1484 1096 1492 1104
rect 1548 1096 1556 1104
rect 1628 1096 1636 1104
rect 1756 1096 1764 1104
rect 1580 1076 1588 1084
rect 1644 1076 1652 1084
rect 1708 1076 1716 1084
rect 1180 996 1188 1004
rect 1244 1056 1252 1064
rect 1356 1056 1364 1064
rect 1246 1006 1254 1014
rect 1260 1006 1268 1014
rect 1274 1006 1282 1014
rect 1484 1056 1492 1064
rect 1500 1056 1508 1064
rect 1660 1056 1668 1064
rect 1708 1056 1716 1064
rect 1436 956 1444 964
rect 1148 936 1156 944
rect 1484 936 1492 944
rect 1116 916 1124 924
rect 1132 896 1140 904
rect 1100 816 1108 824
rect 956 796 964 804
rect 1100 796 1108 804
rect 1068 736 1076 744
rect 940 716 948 724
rect 844 676 852 684
rect 908 676 916 684
rect 556 656 564 664
rect 636 656 644 664
rect 572 636 580 644
rect 588 556 596 564
rect 764 576 772 584
rect 540 536 548 544
rect 556 516 564 524
rect 748 516 756 524
rect 652 496 660 504
rect 684 496 692 504
rect 540 456 548 464
rect 668 456 676 464
rect 636 436 644 444
rect 652 416 660 424
rect 494 406 502 414
rect 508 406 516 414
rect 522 406 530 414
rect 460 336 468 344
rect 428 316 436 324
rect 156 296 164 304
rect 332 296 340 304
rect 364 296 372 304
rect 396 296 404 304
rect 108 176 116 184
rect 172 276 180 284
rect 220 276 228 284
rect 380 276 388 284
rect 204 256 212 264
rect 268 256 276 264
rect 268 176 276 184
rect 60 136 68 144
rect 140 136 148 144
rect 220 136 228 144
rect 140 116 148 124
rect 156 116 164 124
rect 268 116 276 124
rect 12 96 20 104
rect 444 176 452 184
rect 428 136 436 144
rect 460 136 468 144
rect 652 256 660 264
rect 716 256 724 264
rect 812 636 820 644
rect 956 676 964 684
rect 940 656 948 664
rect 892 636 900 644
rect 860 516 868 524
rect 796 476 804 484
rect 828 456 836 464
rect 748 356 756 364
rect 764 316 772 324
rect 764 276 772 284
rect 684 176 692 184
rect 716 156 724 164
rect 764 156 772 164
rect 444 116 452 124
rect 636 116 644 124
rect 572 16 580 24
rect 604 16 612 24
rect 494 6 502 14
rect 508 6 516 14
rect 522 6 530 14
rect 972 596 980 604
rect 924 356 932 364
rect 1116 576 1124 584
rect 1132 576 1140 584
rect 1100 556 1108 564
rect 1132 556 1140 564
rect 1244 916 1252 924
rect 1212 896 1220 904
rect 1452 916 1460 924
rect 1404 856 1412 864
rect 1484 896 1492 904
rect 1468 856 1476 864
rect 1788 1016 1796 1024
rect 1628 956 1636 964
rect 1724 936 1732 944
rect 1548 916 1556 924
rect 1788 956 1796 964
rect 1628 896 1636 904
rect 1212 836 1220 844
rect 1420 836 1428 844
rect 1532 836 1540 844
rect 1196 816 1204 824
rect 1180 696 1188 704
rect 1164 636 1172 644
rect 1164 576 1172 584
rect 1308 736 1316 744
rect 1420 736 1428 744
rect 1596 796 1604 804
rect 1596 776 1604 784
rect 1580 736 1588 744
rect 1404 716 1412 724
rect 1452 716 1460 724
rect 1548 716 1556 724
rect 1228 696 1236 704
rect 1356 696 1364 704
rect 1324 676 1332 684
rect 1372 676 1380 684
rect 1324 656 1332 664
rect 1004 536 1012 544
rect 1196 556 1204 564
rect 1164 536 1172 544
rect 1036 516 1044 524
rect 1084 516 1092 524
rect 1116 516 1124 524
rect 1246 606 1254 614
rect 1260 606 1268 614
rect 1274 606 1282 614
rect 1244 576 1252 584
rect 1132 496 1140 504
rect 1212 496 1220 504
rect 972 476 980 484
rect 972 416 980 424
rect 1116 376 1124 384
rect 1052 336 1060 344
rect 1020 316 1028 324
rect 1068 316 1076 324
rect 1116 316 1124 324
rect 1212 476 1220 484
rect 1196 376 1204 384
rect 1436 676 1444 684
rect 1484 676 1492 684
rect 1644 876 1652 884
rect 1788 856 1796 864
rect 1756 836 1764 844
rect 1724 796 1732 804
rect 1628 736 1636 744
rect 1468 656 1476 664
rect 1596 656 1604 664
rect 1468 576 1476 584
rect 1500 576 1508 584
rect 1388 536 1396 544
rect 1340 516 1348 524
rect 1404 516 1412 524
rect 1564 516 1572 524
rect 1340 476 1348 484
rect 1356 476 1364 484
rect 796 296 804 304
rect 908 296 916 304
rect 1036 296 1044 304
rect 1052 296 1060 304
rect 1132 296 1140 304
rect 1180 296 1188 304
rect 1292 296 1300 304
rect 812 276 820 284
rect 956 276 964 284
rect 1068 276 1076 284
rect 1180 276 1188 284
rect 1212 276 1220 284
rect 1244 276 1252 284
rect 780 136 788 144
rect 892 176 900 184
rect 700 116 708 124
rect 732 116 740 124
rect 844 116 852 124
rect 1068 176 1076 184
rect 972 156 980 164
rect 1116 176 1124 184
rect 1148 176 1156 184
rect 1276 256 1284 264
rect 1246 206 1254 214
rect 1260 206 1268 214
rect 1274 206 1282 214
rect 1292 136 1300 144
rect 956 36 964 44
rect 1004 36 1012 44
rect 940 16 948 24
rect 972 16 980 24
rect 1404 296 1412 304
rect 1356 276 1364 284
rect 1468 276 1476 284
rect 1564 256 1572 264
rect 1356 236 1364 244
rect 1404 236 1412 244
rect 1356 136 1364 144
rect 1324 116 1332 124
rect 1404 116 1412 124
rect 1420 116 1428 124
rect 1452 116 1460 124
rect 1548 116 1556 124
rect 1404 16 1412 24
rect 1436 16 1444 24
rect 1612 516 1620 524
rect 1612 496 1620 504
rect 1772 816 1780 824
rect 1740 576 1748 584
rect 1644 536 1652 544
rect 1740 536 1748 544
rect 1692 496 1700 504
rect 1676 476 1684 484
rect 1628 456 1636 464
rect 1676 456 1684 464
rect 1612 296 1620 304
rect 1628 296 1636 304
rect 1580 236 1588 244
rect 1596 236 1604 244
rect 1596 156 1604 164
rect 1708 236 1716 244
rect 1692 216 1700 224
rect 1788 296 1796 304
rect 1772 216 1780 224
rect 1724 136 1732 144
rect 1756 136 1764 144
rect 1628 116 1636 124
rect 1516 16 1524 24
rect 1564 16 1572 24
<< metal3 >>
rect 1240 1414 1288 1416
rect 1240 1406 1244 1414
rect 1254 1406 1260 1414
rect 1268 1406 1274 1414
rect 1284 1406 1288 1414
rect 1240 1404 1288 1406
rect 852 1397 860 1403
rect 1332 1397 1356 1403
rect 1380 1397 1404 1403
rect 1428 1397 1452 1403
rect 301 1377 748 1383
rect 301 1364 307 1377
rect 212 1357 300 1363
rect 500 1357 620 1363
rect 1108 1357 1132 1363
rect 180 1337 220 1343
rect 228 1337 268 1343
rect 340 1337 396 1343
rect 404 1337 652 1343
rect 749 1337 780 1343
rect 100 1317 124 1323
rect 180 1317 284 1323
rect 340 1317 492 1323
rect 749 1323 755 1337
rect 836 1337 908 1343
rect 1181 1337 1228 1343
rect 612 1317 755 1323
rect 772 1317 860 1323
rect 1181 1323 1187 1337
rect 1028 1317 1187 1323
rect 1204 1317 1276 1323
rect 1316 1317 1468 1323
rect -19 1297 12 1303
rect 132 1297 188 1303
rect 244 1297 348 1303
rect 388 1297 412 1303
rect 740 1297 796 1303
rect 1140 1297 1372 1303
rect 237 1283 243 1296
rect 116 1277 243 1283
rect 292 1277 380 1283
rect 388 1277 620 1283
rect 692 1277 844 1283
rect 488 1214 536 1216
rect 488 1206 492 1214
rect 502 1206 508 1214
rect 516 1206 522 1214
rect 532 1206 536 1214
rect 488 1204 536 1206
rect 836 1197 924 1203
rect 1700 1157 1827 1163
rect 356 1137 428 1143
rect 612 1137 860 1143
rect 68 1117 220 1123
rect 628 1117 700 1123
rect 1460 1117 1660 1123
rect 1796 1117 1827 1123
rect -19 1097 44 1103
rect 52 1097 140 1103
rect 532 1097 604 1103
rect 772 1097 796 1103
rect 852 1097 924 1103
rect 964 1097 1116 1103
rect 1220 1097 1356 1103
rect 1364 1097 1484 1103
rect 1556 1097 1628 1103
rect 1636 1097 1756 1103
rect 132 1077 188 1083
rect 452 1077 588 1083
rect 660 1077 844 1083
rect 868 1077 956 1083
rect 1140 1077 1196 1083
rect 1588 1077 1644 1083
rect 1652 1077 1708 1083
rect 1789 1077 1827 1083
rect -19 1057 3 1063
rect -3 1043 3 1057
rect 36 1057 108 1063
rect 164 1057 396 1063
rect 436 1057 508 1063
rect 724 1057 780 1063
rect 788 1057 908 1063
rect 1252 1057 1356 1063
rect 1364 1057 1484 1063
rect 1508 1057 1660 1063
rect 1789 1063 1795 1077
rect 1716 1057 1795 1063
rect -3 1037 92 1043
rect 109 1043 115 1056
rect 109 1037 188 1043
rect 196 1037 204 1043
rect 260 1017 636 1023
rect 676 1017 716 1023
rect 1796 1017 1827 1023
rect 1240 1014 1288 1016
rect 1240 1006 1244 1014
rect 1254 1006 1260 1014
rect 1268 1006 1274 1014
rect 1284 1006 1288 1014
rect 1240 1004 1288 1006
rect 548 997 972 1003
rect 980 997 1180 1003
rect 340 977 540 983
rect 564 977 924 983
rect 1805 977 1827 983
rect 100 957 396 963
rect 692 957 860 963
rect 1444 957 1628 963
rect 1805 963 1811 977
rect 1796 957 1811 963
rect -19 937 12 943
rect 20 937 60 943
rect 84 937 220 943
rect 260 937 284 943
rect 484 937 860 943
rect 1092 937 1148 943
rect 1156 937 1484 943
rect 1732 937 1740 943
rect 1748 937 1827 943
rect 180 917 204 923
rect 212 917 460 923
rect 676 917 732 923
rect 884 917 908 923
rect 1124 917 1244 923
rect 1252 917 1452 923
rect 1460 917 1548 923
rect -19 897 44 903
rect 52 897 76 903
rect 164 897 236 903
rect 356 897 556 903
rect 628 897 972 903
rect 1060 897 1132 903
rect 1140 897 1212 903
rect 1492 897 1628 903
rect 196 877 380 883
rect 580 877 684 883
rect 1821 883 1827 903
rect 1652 877 1827 883
rect 381 863 387 876
rect 381 857 780 863
rect 1412 857 1468 863
rect 1476 857 1788 863
rect 292 837 860 843
rect 1220 837 1420 843
rect 1540 837 1756 843
rect 1821 843 1827 863
rect 1780 837 1827 843
rect 228 817 444 823
rect 1108 817 1196 823
rect 1780 817 1827 823
rect 488 814 536 816
rect 488 806 492 814
rect 502 806 508 814
rect 516 806 522 814
rect 532 806 536 814
rect 488 804 536 806
rect 580 797 620 803
rect 964 797 1100 803
rect 1108 797 1596 803
rect 1732 797 1772 803
rect 452 777 604 783
rect 644 777 876 783
rect 1604 777 1827 783
rect 612 757 668 763
rect 836 757 892 763
rect -19 737 12 743
rect 84 737 172 743
rect 196 737 252 743
rect 260 737 300 743
rect 596 737 668 743
rect 676 737 844 743
rect 852 737 1068 743
rect 1076 737 1308 743
rect 1316 737 1420 743
rect 1588 737 1628 743
rect 1636 737 1827 743
rect 52 717 60 723
rect 324 717 540 723
rect 548 717 700 723
rect 788 717 796 723
rect 804 717 940 723
rect 1412 717 1452 723
rect 1460 717 1548 723
rect -19 697 92 703
rect 100 697 348 703
rect 596 697 636 703
rect 660 697 684 703
rect 1188 697 1228 703
rect 1236 697 1356 703
rect 1364 697 1827 703
rect 692 677 716 683
rect 740 677 764 683
rect 852 677 908 683
rect 964 677 1004 683
rect 1332 677 1372 683
rect 1444 677 1484 683
rect -19 657 140 663
rect 148 657 556 663
rect 564 657 636 663
rect 948 657 1324 663
rect 1476 657 1596 663
rect 100 637 124 643
rect 420 637 572 643
rect 820 637 892 643
rect 900 637 1164 643
rect 212 617 236 623
rect 244 617 316 623
rect 324 617 412 623
rect 1240 614 1288 616
rect 1240 606 1244 614
rect 1254 606 1260 614
rect 1268 606 1274 614
rect 1284 606 1288 614
rect 1240 604 1288 606
rect -19 577 220 583
rect 308 577 428 583
rect 772 577 1116 583
rect 1172 577 1244 583
rect 1476 577 1500 583
rect 164 557 332 563
rect 372 557 588 563
rect 1108 557 1132 563
rect 1140 557 1196 563
rect -19 537 60 543
rect 228 537 332 543
rect 420 537 540 543
rect 548 537 1004 543
rect 1012 537 1164 543
rect 1396 537 1644 543
rect 1748 537 1827 543
rect 116 517 172 523
rect 324 517 396 523
rect 436 517 556 523
rect 564 517 748 523
rect 868 517 1036 523
rect 1092 517 1116 523
rect 1348 517 1404 523
rect 1412 517 1564 523
rect -19 497 12 503
rect 340 497 444 503
rect 660 497 684 503
rect 1140 497 1212 503
rect 1620 497 1692 503
rect 228 477 796 483
rect 980 477 1212 483
rect 1220 477 1340 483
rect 1348 477 1356 483
rect 1821 483 1827 503
rect 1684 477 1827 483
rect 420 457 540 463
rect 676 457 828 463
rect 1636 457 1676 463
rect 276 437 636 443
rect 644 437 1132 443
rect 660 417 812 423
rect 820 417 972 423
rect 488 414 536 416
rect 488 406 492 414
rect 502 406 508 414
rect 516 406 522 414
rect 532 406 536 414
rect 488 404 536 406
rect 148 377 380 383
rect 388 377 755 383
rect 749 364 755 377
rect 1124 377 1196 383
rect 324 357 412 363
rect 756 357 924 363
rect 356 337 460 343
rect 468 337 1052 343
rect 100 317 252 323
rect 436 317 764 323
rect 1028 317 1068 323
rect 1124 317 1132 323
rect 84 297 156 303
rect 340 297 364 303
rect 404 297 780 303
rect 804 297 908 303
rect 916 297 1036 303
rect 1060 297 1132 303
rect 1188 297 1292 303
rect 1412 297 1612 303
rect 1620 297 1628 303
rect 1796 297 1827 303
rect 180 277 220 283
rect 228 277 380 283
rect 772 277 812 283
rect 964 277 1004 283
rect 1012 277 1068 283
rect 1188 277 1212 283
rect 1220 277 1244 283
rect 1364 277 1468 283
rect 212 257 268 263
rect 660 257 716 263
rect 1284 257 1564 263
rect 980 237 1356 243
rect 1364 237 1404 243
rect 1412 237 1580 243
rect 1588 237 1596 243
rect 1620 237 1708 243
rect 1700 217 1772 223
rect 1240 214 1288 216
rect 1240 206 1244 214
rect 1254 206 1260 214
rect 1268 206 1274 214
rect 1284 206 1288 214
rect 1240 204 1288 206
rect 116 177 268 183
rect 276 177 444 183
rect 452 177 684 183
rect 692 177 892 183
rect 900 177 972 183
rect 1076 177 1107 183
rect 724 157 764 163
rect 772 157 972 163
rect 1101 163 1107 177
rect 1124 177 1148 183
rect 1101 157 1596 163
rect -19 137 60 143
rect 148 137 220 143
rect 436 137 460 143
rect 477 137 780 143
rect 164 117 268 123
rect 276 117 444 123
rect 477 123 483 137
rect 1300 137 1356 143
rect 1732 137 1756 143
rect 452 117 483 123
rect 644 117 700 123
rect 708 117 732 123
rect 820 117 844 123
rect 1332 117 1404 123
rect 1428 117 1452 123
rect 1556 117 1628 123
rect -19 97 12 103
rect 964 37 1004 43
rect 580 17 604 23
rect 948 17 972 23
rect 1412 17 1436 23
rect 1524 17 1564 23
rect 488 14 536 16
rect 488 6 492 14
rect 502 6 508 14
rect 516 6 522 14
rect 532 6 536 14
rect 488 4 536 6
<< m4contact >>
rect 1244 1406 1246 1414
rect 1246 1406 1252 1414
rect 1260 1406 1268 1414
rect 1276 1406 1282 1414
rect 1282 1406 1284 1414
rect 844 1396 852 1404
rect 492 1206 494 1214
rect 494 1206 500 1214
rect 508 1206 516 1214
rect 524 1206 530 1214
rect 530 1206 532 1214
rect 844 1096 852 1104
rect 1244 1006 1246 1014
rect 1246 1006 1252 1014
rect 1260 1006 1268 1014
rect 1276 1006 1282 1014
rect 1282 1006 1284 1014
rect 972 996 980 1004
rect 44 956 52 964
rect 1740 936 1748 944
rect 1772 836 1780 844
rect 492 806 494 814
rect 494 806 500 814
rect 508 806 516 814
rect 524 806 530 814
rect 530 806 532 814
rect 1772 796 1780 804
rect 44 716 52 724
rect 780 716 788 724
rect 268 676 276 684
rect 1004 676 1012 684
rect 1244 606 1246 614
rect 1246 606 1252 614
rect 1260 606 1268 614
rect 1276 606 1282 614
rect 1282 606 1284 614
rect 972 596 980 604
rect 1132 576 1140 584
rect 1740 576 1748 584
rect 1612 516 1620 524
rect 268 436 276 444
rect 1132 436 1140 444
rect 812 416 820 424
rect 492 406 494 414
rect 494 406 500 414
rect 508 406 516 414
rect 524 406 530 414
rect 530 406 532 414
rect 140 376 148 384
rect 1132 316 1140 324
rect 780 296 788 304
rect 1004 276 1012 284
rect 972 236 980 244
rect 1612 236 1620 244
rect 1244 206 1246 214
rect 1246 206 1252 214
rect 1260 206 1268 214
rect 1276 206 1282 214
rect 1282 206 1284 214
rect 972 176 980 184
rect 140 116 148 124
rect 812 116 820 124
rect 492 6 494 14
rect 494 6 500 14
rect 508 6 516 14
rect 524 6 530 14
rect 530 6 532 14
<< metal4 >>
rect 488 1214 536 1440
rect 1240 1414 1288 1440
rect 1240 1406 1244 1414
rect 1252 1406 1260 1414
rect 1268 1406 1276 1414
rect 1284 1406 1288 1414
rect 488 1206 492 1214
rect 500 1206 508 1214
rect 516 1206 524 1214
rect 532 1206 536 1214
rect 42 964 54 966
rect 42 956 44 964
rect 52 956 54 964
rect 42 724 54 956
rect 42 716 44 724
rect 52 716 54 724
rect 42 714 54 716
rect 488 814 536 1206
rect 842 1404 854 1406
rect 842 1396 844 1404
rect 852 1396 854 1404
rect 842 1104 854 1396
rect 842 1096 844 1104
rect 852 1096 854 1104
rect 842 1094 854 1096
rect 1240 1014 1288 1406
rect 1240 1006 1244 1014
rect 1252 1006 1260 1014
rect 1268 1006 1276 1014
rect 1284 1006 1288 1014
rect 488 806 492 814
rect 500 806 508 814
rect 516 806 524 814
rect 532 806 536 814
rect 266 684 278 686
rect 266 676 268 684
rect 276 676 278 684
rect 266 444 278 676
rect 266 436 268 444
rect 276 436 278 444
rect 266 434 278 436
rect 488 414 536 806
rect 970 1004 982 1006
rect 970 996 972 1004
rect 980 996 982 1004
rect 488 406 492 414
rect 500 406 508 414
rect 516 406 524 414
rect 532 406 536 414
rect 138 384 150 386
rect 138 376 140 384
rect 148 376 150 384
rect 138 124 150 376
rect 138 116 140 124
rect 148 116 150 124
rect 138 114 150 116
rect 488 14 536 406
rect 778 724 790 726
rect 778 716 780 724
rect 788 716 790 724
rect 778 304 790 716
rect 970 604 982 996
rect 970 596 972 604
rect 980 596 982 604
rect 778 296 780 304
rect 788 296 790 304
rect 778 294 790 296
rect 810 424 822 426
rect 810 416 812 424
rect 820 416 822 424
rect 810 124 822 416
rect 970 244 982 596
rect 1002 684 1014 686
rect 1002 676 1004 684
rect 1012 676 1014 684
rect 1002 284 1014 676
rect 1240 614 1288 1006
rect 1240 606 1244 614
rect 1252 606 1260 614
rect 1268 606 1276 614
rect 1284 606 1288 614
rect 1130 584 1142 586
rect 1130 576 1132 584
rect 1140 576 1142 584
rect 1130 444 1142 576
rect 1130 436 1132 444
rect 1140 436 1142 444
rect 1130 324 1142 436
rect 1130 316 1132 324
rect 1140 316 1142 324
rect 1130 314 1142 316
rect 1002 276 1004 284
rect 1012 276 1014 284
rect 1002 274 1014 276
rect 970 236 972 244
rect 980 236 982 244
rect 970 184 982 236
rect 970 176 972 184
rect 980 176 982 184
rect 970 174 982 176
rect 1240 214 1288 606
rect 1738 944 1750 946
rect 1738 936 1740 944
rect 1748 936 1750 944
rect 1738 584 1750 936
rect 1770 844 1782 846
rect 1770 836 1772 844
rect 1780 836 1782 844
rect 1770 804 1782 836
rect 1770 796 1772 804
rect 1780 796 1782 804
rect 1770 794 1782 796
rect 1738 576 1740 584
rect 1748 576 1750 584
rect 1738 574 1750 576
rect 1610 524 1622 526
rect 1610 516 1612 524
rect 1620 516 1622 524
rect 1610 244 1622 516
rect 1610 236 1612 244
rect 1620 236 1622 244
rect 1610 234 1622 236
rect 1240 206 1244 214
rect 1252 206 1260 214
rect 1268 206 1276 214
rect 1284 206 1288 214
rect 810 116 812 124
rect 820 116 822 124
rect 810 114 822 116
rect 488 6 492 14
rect 500 6 508 14
rect 516 6 524 14
rect 532 6 536 14
rect 488 -40 536 6
rect 1240 -40 1288 206
use BUFX2  BUFX2_21
timestamp 1651685240
transform -1 0 56 0 -1 210
box -4 -6 52 206
use BUFX2  BUFX2_25
timestamp 1651685240
transform -1 0 104 0 -1 210
box -4 -6 52 206
use AND2X2  AND2X2_10
timestamp 1651685240
transform -1 0 168 0 -1 210
box -4 -6 68 206
use NOR3X1  NOR3X1_16
timestamp 1651685240
transform -1 0 136 0 1 210
box -4 -6 132 206
use OR2X2  OR2X2_3
timestamp 1651685240
transform -1 0 200 0 1 210
box -4 -6 68 206
use BUFX2  BUFX2_22
timestamp 1651685240
transform -1 0 216 0 -1 210
box -4 -6 52 206
use NOR3X1  NOR3X1_17
timestamp 1651685240
transform 1 0 216 0 -1 210
box -4 -6 132 206
use OAI21X1  OAI21X1_5
timestamp 1651685240
transform 1 0 200 0 1 210
box -4 -6 68 206
use INVX1  INVX1_10
timestamp 1651685240
transform -1 0 296 0 1 210
box -4 -6 36 206
use BUFX2  BUFX2_20
timestamp 1651685240
transform -1 0 392 0 -1 210
box -4 -6 52 206
use NOR3X1  NOR3X1_15
timestamp 1651685240
transform 1 0 392 0 -1 210
box -4 -6 132 206
use NAND3X1  NAND3X1_6
timestamp 1651685240
transform -1 0 360 0 1 210
box -4 -6 68 206
use AOI21X1  AOI21X1_4
timestamp 1651685240
transform -1 0 424 0 1 210
box -4 -6 68 206
use FILL  FILL_0_0_0
timestamp 1651685240
transform 1 0 520 0 -1 210
box -4 -6 20 206
use FILL  FILL_0_0_1
timestamp 1651685240
transform 1 0 536 0 -1 210
box -4 -6 20 206
use FILL  FILL_0_0_2
timestamp 1651685240
transform 1 0 552 0 -1 210
box -4 -6 20 206
use XNOR2X1  XNOR2X1_8
timestamp 1651685240
transform 1 0 424 0 1 210
box -4 -6 116 206
use FILL  FILL_1_0_0
timestamp 1651685240
transform -1 0 552 0 1 210
box -4 -6 20 206
use FILL  FILL_1_0_1
timestamp 1651685240
transform -1 0 568 0 1 210
box -4 -6 20 206
use BUFX2  BUFX2_23
timestamp 1651685240
transform 1 0 568 0 -1 210
box -4 -6 52 206
use NOR2X1  NOR2X1_9
timestamp 1651685240
transform -1 0 664 0 -1 210
box -4 -6 52 206
use AND2X2  AND2X2_4
timestamp 1651685240
transform -1 0 728 0 -1 210
box -4 -6 68 206
use FILL  FILL_1_0_2
timestamp 1651685240
transform -1 0 584 0 1 210
box -4 -6 20 206
use NOR3X1  NOR3X1_18
timestamp 1651685240
transform -1 0 712 0 1 210
box -4 -6 132 206
use NAND2X1  NAND2X1_4
timestamp 1651685240
transform -1 0 776 0 -1 210
box -4 -6 52 206
use NOR3X1  NOR3X1_14
timestamp 1651685240
transform -1 0 904 0 -1 210
box -4 -6 132 206
use INVX1  INVX1_12
timestamp 1651685240
transform 1 0 712 0 1 210
box -4 -6 36 206
use OAI21X1  OAI21X1_17
timestamp 1651685240
transform 1 0 744 0 1 210
box -4 -6 68 206
use XNOR2X1  XNOR2X1_7
timestamp 1651685240
transform -1 0 920 0 1 210
box -4 -6 116 206
use BUFX2  BUFX2_19
timestamp 1651685240
transform 1 0 904 0 -1 210
box -4 -6 52 206
use NOR2X1  NOR2X1_8
timestamp 1651685240
transform 1 0 952 0 -1 210
box -4 -6 52 206
use BUFX2  BUFX2_17
timestamp 1651685240
transform -1 0 968 0 1 210
box -4 -6 52 206
use XOR2X1  XOR2X1_8
timestamp 1651685240
transform -1 0 1112 0 -1 210
box -4 -6 116 206
use INVX1  INVX1_13
timestamp 1651685240
transform 1 0 968 0 1 210
box -4 -6 36 206
use OAI21X1  OAI21X1_16
timestamp 1651685240
transform 1 0 1000 0 1 210
box -4 -6 68 206
use OAI21X1  OAI21X1_15
timestamp 1651685240
transform 1 0 1064 0 1 210
box -4 -6 68 206
use XOR2X1  XOR2X1_5
timestamp 1651685240
transform 1 0 1112 0 -1 210
box -4 -6 116 206
use FILL  FILL_0_1_0
timestamp 1651685240
transform -1 0 1240 0 -1 210
box -4 -6 20 206
use NAND2X1  NAND2X1_19
timestamp 1651685240
transform 1 0 1128 0 1 210
box -4 -6 52 206
use NOR2X1  NOR2X1_7
timestamp 1651685240
transform 1 0 1176 0 1 210
box -4 -6 52 206
use FILL  FILL_1_1_0
timestamp 1651685240
transform 1 0 1224 0 1 210
box -4 -6 20 206
use FILL  FILL_0_1_1
timestamp 1651685240
transform -1 0 1256 0 -1 210
box -4 -6 20 206
use FILL  FILL_0_1_2
timestamp 1651685240
transform -1 0 1272 0 -1 210
box -4 -6 20 206
use NOR3X1  NOR3X1_10
timestamp 1651685240
transform -1 0 1400 0 -1 210
box -4 -6 132 206
use FILL  FILL_1_1_1
timestamp 1651685240
transform 1 0 1240 0 1 210
box -4 -6 20 206
use FILL  FILL_1_1_2
timestamp 1651685240
transform 1 0 1256 0 1 210
box -4 -6 20 206
use OAI21X1  OAI21X1_13
timestamp 1651685240
transform 1 0 1272 0 1 210
box -4 -6 68 206
use NOR3X1  NOR3X1_6
timestamp 1651685240
transform -1 0 1464 0 1 210
box -4 -6 132 206
use BUFX2  BUFX2_15
timestamp 1651685240
transform 1 0 1400 0 -1 210
box -4 -6 52 206
use BUFX2  BUFX2_11
timestamp 1651685240
transform 1 0 1448 0 -1 210
box -4 -6 52 206
use NOR3X1  NOR3X1_13
timestamp 1651685240
transform -1 0 1624 0 -1 210
box -4 -6 132 206
use XOR2X1  XOR2X1_6
timestamp 1651685240
transform 1 0 1464 0 1 210
box -4 -6 116 206
use BUFX2  BUFX2_18
timestamp 1651685240
transform 1 0 1624 0 -1 210
box -4 -6 52 206
use NOR3X1  NOR3X1_11
timestamp 1651685240
transform 1 0 1576 0 1 210
box -4 -6 132 206
use AND2X2  AND2X2_2
timestamp 1651685240
transform -1 0 1736 0 -1 210
box -4 -6 68 206
use BUFX2  BUFX2_16
timestamp 1651685240
transform -1 0 1784 0 -1 210
box -4 -6 52 206
use BUFX2  BUFX2_29
timestamp 1651685240
transform 1 0 1704 0 1 210
box -4 -6 52 206
use FILL  FILL_2_1
timestamp 1651685240
transform 1 0 1752 0 1 210
box -4 -6 20 206
use FILL  FILL_2_2
timestamp 1651685240
transform 1 0 1768 0 1 210
box -4 -6 20 206
use FILL  FILL_1_1
timestamp 1651685240
transform -1 0 1800 0 -1 210
box -4 -6 20 206
use FILL  FILL_2_3
timestamp 1651685240
transform 1 0 1784 0 1 210
box -4 -6 20 206
use BUFX2  BUFX2_31
timestamp 1651685240
transform -1 0 56 0 -1 610
box -4 -6 52 206
use BUFX2  BUFX2_32
timestamp 1651685240
transform -1 0 104 0 -1 610
box -4 -6 52 206
use NAND2X1  NAND2X1_5
timestamp 1651685240
transform -1 0 152 0 -1 610
box -4 -6 52 206
use AND2X2  AND2X2_5
timestamp 1651685240
transform 1 0 152 0 -1 610
box -4 -6 68 206
use XNOR2X1  XNOR2X1_1
timestamp 1651685240
transform -1 0 328 0 -1 610
box -4 -6 116 206
use NOR2X1  NOR2X1_11
timestamp 1651685240
transform -1 0 376 0 -1 610
box -4 -6 52 206
use AOI21X1  AOI21X1_5
timestamp 1651685240
transform -1 0 440 0 -1 610
box -4 -6 68 206
use INVX1  INVX1_9
timestamp 1651685240
transform 1 0 440 0 -1 610
box -4 -6 36 206
use FILL  FILL_2_0_0
timestamp 1651685240
transform 1 0 472 0 -1 610
box -4 -6 20 206
use FILL  FILL_2_0_1
timestamp 1651685240
transform 1 0 488 0 -1 610
box -4 -6 20 206
use FILL  FILL_2_0_2
timestamp 1651685240
transform 1 0 504 0 -1 610
box -4 -6 20 206
use NAND3X1  NAND3X1_5
timestamp 1651685240
transform 1 0 520 0 -1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_4
timestamp 1651685240
transform 1 0 584 0 -1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_13
timestamp 1651685240
transform 1 0 648 0 -1 610
box -4 -6 52 206
use INVX1  INVX1_14
timestamp 1651685240
transform -1 0 728 0 -1 610
box -4 -6 36 206
use NOR2X1  NOR2X1_10
timestamp 1651685240
transform -1 0 776 0 -1 610
box -4 -6 52 206
use BUFX2  BUFX2_3
timestamp 1651685240
transform -1 0 824 0 -1 610
box -4 -6 52 206
use NAND2X1  NAND2X1_10
timestamp 1651685240
transform -1 0 872 0 -1 610
box -4 -6 52 206
use NOR3X1  NOR3X1_12
timestamp 1651685240
transform -1 0 1000 0 -1 610
box -4 -6 132 206
use NAND2X1  NAND2X1_20
timestamp 1651685240
transform -1 0 1048 0 -1 610
box -4 -6 52 206
use AND2X2  AND2X2_3
timestamp 1651685240
transform -1 0 1112 0 -1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_3
timestamp 1651685240
transform -1 0 1160 0 -1 610
box -4 -6 52 206
use NAND2X1  NAND2X1_18
timestamp 1651685240
transform -1 0 1208 0 -1 610
box -4 -6 52 206
use BUFX2  BUFX2_1
timestamp 1651685240
transform -1 0 1256 0 -1 610
box -4 -6 52 206
use FILL  FILL_2_1_0
timestamp 1651685240
transform 1 0 1256 0 -1 610
box -4 -6 20 206
use FILL  FILL_2_1_1
timestamp 1651685240
transform 1 0 1272 0 -1 610
box -4 -6 20 206
use FILL  FILL_2_1_2
timestamp 1651685240
transform 1 0 1288 0 -1 610
box -4 -6 20 206
use BUFX2  BUFX2_4
timestamp 1651685240
transform 1 0 1304 0 -1 610
box -4 -6 52 206
use NOR2X1  NOR2X1_21
timestamp 1651685240
transform -1 0 1400 0 -1 610
box -4 -6 52 206
use XOR2X1  XOR2X1_3
timestamp 1651685240
transform 1 0 1400 0 -1 610
box -4 -6 116 206
use NOR3X1  NOR3X1_7
timestamp 1651685240
transform 1 0 1512 0 -1 610
box -4 -6 132 206
use BUFX2  BUFX2_24
timestamp 1651685240
transform 1 0 1640 0 -1 610
box -4 -6 52 206
use BUFX2  BUFX2_12
timestamp 1651685240
transform 1 0 1688 0 -1 610
box -4 -6 52 206
use NOR2X1  NOR2X1_3
timestamp 1651685240
transform 1 0 1736 0 -1 610
box -4 -6 52 206
use FILL  FILL_3_1
timestamp 1651685240
transform -1 0 1800 0 -1 610
box -4 -6 20 206
use BUFX2  BUFX2_36
timestamp 1651685240
transform -1 0 56 0 1 610
box -4 -6 52 206
use NOR2X1  NOR2X1_15
timestamp 1651685240
transform -1 0 104 0 1 610
box -4 -6 52 206
use NOR2X1  NOR2X1_12
timestamp 1651685240
transform -1 0 152 0 1 610
box -4 -6 52 206
use NAND3X1  NAND3X1_1
timestamp 1651685240
transform -1 0 216 0 1 610
box -4 -6 68 206
use NAND3X1  NAND3X1_8
timestamp 1651685240
transform 1 0 216 0 1 610
box -4 -6 68 206
use NAND3X1  NAND3X1_3
timestamp 1651685240
transform -1 0 344 0 1 610
box -4 -6 68 206
use XNOR2X1  XNOR2X1_2
timestamp 1651685240
transform -1 0 456 0 1 610
box -4 -6 116 206
use FILL  FILL_3_0_0
timestamp 1651685240
transform -1 0 472 0 1 610
box -4 -6 20 206
use FILL  FILL_3_0_1
timestamp 1651685240
transform -1 0 488 0 1 610
box -4 -6 20 206
use FILL  FILL_3_0_2
timestamp 1651685240
transform -1 0 504 0 1 610
box -4 -6 20 206
use OAI21X1  OAI21X1_8
timestamp 1651685240
transform -1 0 568 0 1 610
box -4 -6 68 206
use AOI21X1  AOI21X1_6
timestamp 1651685240
transform -1 0 632 0 1 610
box -4 -6 68 206
use INVX1  INVX1_8
timestamp 1651685240
transform 1 0 632 0 1 610
box -4 -6 36 206
use NAND3X1  NAND3X1_4
timestamp 1651685240
transform 1 0 664 0 1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_14
timestamp 1651685240
transform -1 0 776 0 1 610
box -4 -6 52 206
use AOI22X1  AOI22X1_2
timestamp 1651685240
transform 1 0 776 0 1 610
box -4 -6 84 206
use NAND3X1  NAND3X1_10
timestamp 1651685240
transform 1 0 856 0 1 610
box -4 -6 68 206
use INVX1  INVX1_1
timestamp 1651685240
transform -1 0 952 0 1 610
box -4 -6 36 206
use XOR2X1  XOR2X1_7
timestamp 1651685240
transform -1 0 1064 0 1 610
box -4 -6 116 206
use OAI21X1  OAI21X1_14
timestamp 1651685240
transform -1 0 1128 0 1 610
box -4 -6 68 206
use BUFX2  BUFX2_7
timestamp 1651685240
transform -1 0 1176 0 1 610
box -4 -6 52 206
use BUFX2  BUFX2_8
timestamp 1651685240
transform 1 0 1176 0 1 610
box -4 -6 52 206
use BUFX2  BUFX2_6
timestamp 1651685240
transform 1 0 1224 0 1 610
box -4 -6 52 206
use FILL  FILL_3_1_0
timestamp 1651685240
transform -1 0 1288 0 1 610
box -4 -6 20 206
use FILL  FILL_3_1_1
timestamp 1651685240
transform -1 0 1304 0 1 610
box -4 -6 20 206
use FILL  FILL_3_1_2
timestamp 1651685240
transform -1 0 1320 0 1 610
box -4 -6 20 206
use BUFX2  BUFX2_5
timestamp 1651685240
transform -1 0 1368 0 1 610
box -4 -6 52 206
use NAND2X1  NAND2X1_17
timestamp 1651685240
transform 1 0 1368 0 1 610
box -4 -6 52 206
use OAI21X1  OAI21X1_10
timestamp 1651685240
transform -1 0 1480 0 1 610
box -4 -6 68 206
use XOR2X1  XOR2X1_4
timestamp 1651685240
transform 1 0 1480 0 1 610
box -4 -6 116 206
use NOR2X1  NOR2X1_4
timestamp 1651685240
transform 1 0 1592 0 1 610
box -4 -6 52 206
use BUFX2  BUFX2_30
timestamp 1651685240
transform -1 0 1688 0 1 610
box -4 -6 52 206
use BUFX2  BUFX2_35
timestamp 1651685240
transform 1 0 1688 0 1 610
box -4 -6 52 206
use BUFX2  BUFX2_33
timestamp 1651685240
transform 1 0 1736 0 1 610
box -4 -6 52 206
use FILL  FILL_4_1
timestamp 1651685240
transform 1 0 1784 0 1 610
box -4 -6 20 206
use NOR2X1  NOR2X1_13
timestamp 1651685240
transform 1 0 8 0 -1 1010
box -4 -6 52 206
use AND2X2  AND2X2_8
timestamp 1651685240
transform 1 0 56 0 -1 1010
box -4 -6 68 206
use MUX2X1  MUX2X1_1
timestamp 1651685240
transform -1 0 216 0 -1 1010
box -4 -6 100 206
use OAI21X1  OAI21X1_7
timestamp 1651685240
transform 1 0 216 0 -1 1010
box -4 -6 68 206
use XNOR2X1  XNOR2X1_4
timestamp 1651685240
transform 1 0 280 0 -1 1010
box -4 -6 116 206
use INVX1  INVX1_5
timestamp 1651685240
transform 1 0 392 0 -1 1010
box -4 -6 36 206
use NAND3X1  NAND3X1_2
timestamp 1651685240
transform 1 0 424 0 -1 1010
box -4 -6 68 206
use FILL  FILL_4_0_0
timestamp 1651685240
transform -1 0 504 0 -1 1010
box -4 -6 20 206
use FILL  FILL_4_0_1
timestamp 1651685240
transform -1 0 520 0 -1 1010
box -4 -6 20 206
use FILL  FILL_4_0_2
timestamp 1651685240
transform -1 0 536 0 -1 1010
box -4 -6 20 206
use NAND3X1  NAND3X1_9
timestamp 1651685240
transform -1 0 600 0 -1 1010
box -4 -6 68 206
use NAND2X1  NAND2X1_11
timestamp 1651685240
transform 1 0 600 0 -1 1010
box -4 -6 52 206
use NAND3X1  NAND3X1_7
timestamp 1651685240
transform 1 0 648 0 -1 1010
box -4 -6 68 206
use NOR3X1  NOR3X1_1
timestamp 1651685240
transform -1 0 840 0 -1 1010
box -4 -6 132 206
use INVX1  INVX1_3
timestamp 1651685240
transform -1 0 872 0 -1 1010
box -4 -6 36 206
use NOR2X1  NOR2X1_19
timestamp 1651685240
transform -1 0 920 0 -1 1010
box -4 -6 52 206
use NOR3X1  NOR3X1_2
timestamp 1651685240
transform 1 0 920 0 -1 1010
box -4 -6 132 206
use OAI21X1  OAI21X1_11
timestamp 1651685240
transform -1 0 1112 0 -1 1010
box -4 -6 68 206
use NOR2X1  NOR2X1_5
timestamp 1651685240
transform 1 0 1112 0 -1 1010
box -4 -6 52 206
use BUFX2  BUFX2_2
timestamp 1651685240
transform 1 0 1160 0 -1 1010
box -4 -6 52 206
use NAND2X1  NAND2X1_15
timestamp 1651685240
transform 1 0 1208 0 -1 1010
box -4 -6 52 206
use FILL  FILL_4_1_0
timestamp 1651685240
transform 1 0 1256 0 -1 1010
box -4 -6 20 206
use FILL  FILL_4_1_1
timestamp 1651685240
transform 1 0 1272 0 -1 1010
box -4 -6 20 206
use FILL  FILL_4_1_2
timestamp 1651685240
transform 1 0 1288 0 -1 1010
box -4 -6 20 206
use XOR2X1  XOR2X1_1
timestamp 1651685240
transform 1 0 1304 0 -1 1010
box -4 -6 116 206
use OAI21X1  OAI21X1_9
timestamp 1651685240
transform -1 0 1480 0 -1 1010
box -4 -6 68 206
use NAND2X1  NAND2X1_2
timestamp 1651685240
transform -1 0 1528 0 -1 1010
box -4 -6 52 206
use NAND2X1  NAND2X1_16
timestamp 1651685240
transform 1 0 1528 0 -1 1010
box -4 -6 52 206
use NAND2X1  NAND2X1_9
timestamp 1651685240
transform 1 0 1576 0 -1 1010
box -4 -6 52 206
use XOR2X1  XOR2X1_2
timestamp 1651685240
transform 1 0 1624 0 -1 1010
box -4 -6 116 206
use BUFX2  BUFX2_26
timestamp 1651685240
transform 1 0 1736 0 -1 1010
box -4 -6 52 206
use FILL  FILL_5_1
timestamp 1651685240
transform -1 0 1800 0 -1 1010
box -4 -6 20 206
use NAND2X1  NAND2X1_6
timestamp 1651685240
transform 1 0 8 0 1 1010
box -4 -6 52 206
use NOR2X1  NOR2X1_14
timestamp 1651685240
transform -1 0 104 0 1 1010
box -4 -6 52 206
use INVX1  INVX1_4
timestamp 1651685240
transform 1 0 104 0 1 1010
box -4 -6 36 206
use OAI21X1  OAI21X1_2
timestamp 1651685240
transform -1 0 200 0 1 1010
box -4 -6 68 206
use AND2X2  AND2X2_6
timestamp 1651685240
transform 1 0 200 0 1 1010
box -4 -6 68 206
use XNOR2X1  XNOR2X1_3
timestamp 1651685240
transform -1 0 376 0 1 1010
box -4 -6 116 206
use AOI22X1  AOI22X1_1
timestamp 1651685240
transform 1 0 376 0 1 1010
box -4 -6 84 206
use FILL  FILL_5_0_0
timestamp 1651685240
transform 1 0 456 0 1 1010
box -4 -6 20 206
use FILL  FILL_5_0_1
timestamp 1651685240
transform 1 0 472 0 1 1010
box -4 -6 20 206
use FILL  FILL_5_0_2
timestamp 1651685240
transform 1 0 488 0 1 1010
box -4 -6 20 206
use AOI21X1  AOI21X1_1
timestamp 1651685240
transform 1 0 504 0 1 1010
box -4 -6 68 206
use NAND2X1  NAND2X1_12
timestamp 1651685240
transform 1 0 568 0 1 1010
box -4 -6 52 206
use OAI21X1  OAI21X1_1
timestamp 1651685240
transform -1 0 680 0 1 1010
box -4 -6 68 206
use NAND2X1  NAND2X1_8
timestamp 1651685240
transform -1 0 728 0 1 1010
box -4 -6 52 206
use AND2X2  AND2X2_9
timestamp 1651685240
transform -1 0 792 0 1 1010
box -4 -6 68 206
use NOR2X1  NOR2X1_20
timestamp 1651685240
transform 1 0 792 0 1 1010
box -4 -6 52 206
use NAND2X1  NAND2X1_7
timestamp 1651685240
transform -1 0 888 0 1 1010
box -4 -6 52 206
use NOR2X1  NOR2X1_18
timestamp 1651685240
transform 1 0 888 0 1 1010
box -4 -6 52 206
use OAI21X1  OAI21X1_12
timestamp 1651685240
transform 1 0 936 0 1 1010
box -4 -6 68 206
use XNOR2X1  XNOR2X1_5
timestamp 1651685240
transform 1 0 1000 0 1 1010
box -4 -6 116 206
use NOR3X1  NOR3X1_8
timestamp 1651685240
transform -1 0 1240 0 1 1010
box -4 -6 132 206
use FILL  FILL_5_1_0
timestamp 1651685240
transform -1 0 1256 0 1 1010
box -4 -6 20 206
use FILL  FILL_5_1_1
timestamp 1651685240
transform -1 0 1272 0 1 1010
box -4 -6 20 206
use FILL  FILL_5_1_2
timestamp 1651685240
transform -1 0 1288 0 1 1010
box -4 -6 20 206
use NOR3X1  NOR3X1_4
timestamp 1651685240
transform -1 0 1416 0 1 1010
box -4 -6 132 206
use NOR3X1  NOR3X1_5
timestamp 1651685240
transform -1 0 1544 0 1 1010
box -4 -6 132 206
use NAND2X1  NAND2X1_1
timestamp 1651685240
transform -1 0 1592 0 1 1010
box -4 -6 52 206
use AND2X2  AND2X2_1
timestamp 1651685240
transform -1 0 1656 0 1 1010
box -4 -6 68 206
use BUFX2  BUFX2_10
timestamp 1651685240
transform 1 0 1656 0 1 1010
box -4 -6 52 206
use NOR2X1  NOR2X1_1
timestamp 1651685240
transform 1 0 1704 0 1 1010
box -4 -6 52 206
use FILL  FILL_6_1
timestamp 1651685240
transform 1 0 1752 0 1 1010
box -4 -6 20 206
use FILL  FILL_6_2
timestamp 1651685240
transform 1 0 1768 0 1 1010
box -4 -6 20 206
use FILL  FILL_6_3
timestamp 1651685240
transform 1 0 1784 0 1 1010
box -4 -6 20 206
use BUFX2  BUFX2_28
timestamp 1651685240
transform -1 0 56 0 -1 1410
box -4 -6 52 206
use AND2X2  AND2X2_7
timestamp 1651685240
transform -1 0 120 0 -1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_6
timestamp 1651685240
transform -1 0 184 0 -1 1410
box -4 -6 68 206
use NOR2X1  NOR2X1_16
timestamp 1651685240
transform -1 0 232 0 -1 1410
box -4 -6 52 206
use OR2X2  OR2X2_2
timestamp 1651685240
transform -1 0 296 0 -1 1410
box -4 -6 68 206
use INVX1  INVX1_2
timestamp 1651685240
transform 1 0 296 0 -1 1410
box -4 -6 36 206
use OAI21X1  OAI21X1_3
timestamp 1651685240
transform 1 0 328 0 -1 1410
box -4 -6 68 206
use OR2X2  OR2X2_1
timestamp 1651685240
transform 1 0 392 0 -1 1410
box -4 -6 68 206
use NOR2X1  NOR2X1_17
timestamp 1651685240
transform 1 0 456 0 -1 1410
box -4 -6 52 206
use FILL  FILL_6_0_0
timestamp 1651685240
transform -1 0 520 0 -1 1410
box -4 -6 20 206
use FILL  FILL_6_0_1
timestamp 1651685240
transform -1 0 536 0 -1 1410
box -4 -6 20 206
use FILL  FILL_6_0_2
timestamp 1651685240
transform -1 0 552 0 -1 1410
box -4 -6 20 206
use NOR3X1  NOR3X1_3
timestamp 1651685240
transform -1 0 680 0 -1 1410
box -4 -6 132 206
use INVX1  INVX1_6
timestamp 1651685240
transform 1 0 680 0 -1 1410
box -4 -6 36 206
use AOI21X1  AOI21X1_2
timestamp 1651685240
transform -1 0 776 0 -1 1410
box -4 -6 68 206
use OAI22X1  OAI22X1_1
timestamp 1651685240
transform 1 0 776 0 -1 1410
box -4 -6 84 206
use AOI21X1  AOI21X1_3
timestamp 1651685240
transform 1 0 856 0 -1 1410
box -4 -6 68 206
use INVX1  INVX1_7
timestamp 1651685240
transform -1 0 952 0 -1 1410
box -4 -6 36 206
use XNOR2X1  XNOR2X1_6
timestamp 1651685240
transform 1 0 952 0 -1 1410
box -4 -6 116 206
use NOR2X1  NOR2X1_6
timestamp 1651685240
transform -1 0 1112 0 -1 1410
box -4 -6 52 206
use INVX1  INVX1_11
timestamp 1651685240
transform -1 0 1144 0 -1 1410
box -4 -6 36 206
use NOR3X1  NOR3X1_9
timestamp 1651685240
transform -1 0 1272 0 -1 1410
box -4 -6 132 206
use FILL  FILL_6_1_0
timestamp 1651685240
transform 1 0 1272 0 -1 1410
box -4 -6 20 206
use FILL  FILL_6_1_1
timestamp 1651685240
transform 1 0 1288 0 -1 1410
box -4 -6 20 206
use FILL  FILL_6_1_2
timestamp 1651685240
transform 1 0 1304 0 -1 1410
box -4 -6 20 206
use BUFX2  BUFX2_14
timestamp 1651685240
transform 1 0 1320 0 -1 1410
box -4 -6 52 206
use BUFX2  BUFX2_13
timestamp 1651685240
transform 1 0 1368 0 -1 1410
box -4 -6 52 206
use BUFX2  BUFX2_39
timestamp 1651685240
transform 1 0 1416 0 -1 1410
box -4 -6 52 206
use BUFX2  BUFX2_9
timestamp 1651685240
transform 1 0 1464 0 -1 1410
box -4 -6 52 206
use BUFX2  BUFX2_34
timestamp 1651685240
transform 1 0 1512 0 -1 1410
box -4 -6 52 206
use BUFX2  BUFX2_27
timestamp 1651685240
transform 1 0 1560 0 -1 1410
box -4 -6 52 206
use BUFX2  BUFX2_37
timestamp 1651685240
transform 1 0 1608 0 -1 1410
box -4 -6 52 206
use BUFX2  BUFX2_40
timestamp 1651685240
transform 1 0 1656 0 -1 1410
box -4 -6 52 206
use BUFX2  BUFX2_38
timestamp 1651685240
transform 1 0 1704 0 -1 1410
box -4 -6 52 206
use NOR2X1  NOR2X1_2
timestamp 1651685240
transform -1 0 1800 0 -1 1410
box -4 -6 52 206
<< labels >>
flabel metal4 s 488 -40 536 -16 7 FreeSans 24 270 0 0 vdd
port 0 nsew
flabel metal4 s 1240 -40 1288 -16 7 FreeSans 24 270 0 0 gnd
port 1 nsew
flabel metal3 s 1821 1077 1827 1083 3 FreeSans 24 0 0 0 Y[0]
port 2 nsew
flabel metal2 s 1805 1437 1811 1443 3 FreeSans 24 90 0 0 Y[1]
port 3 nsew
flabel metal2 s 1773 1437 1779 1443 3 FreeSans 24 90 0 0 Y[2]
port 4 nsew
flabel metal3 s 1821 1117 1827 1123 3 FreeSans 24 0 0 0 Y[3]
port 5 nsew
flabel metal3 s 1821 977 1827 983 3 FreeSans 24 0 0 0 Y[4]
port 6 nsew
flabel metal3 s 1821 937 1827 943 3 FreeSans 24 0 0 0 Y[5]
port 7 nsew
flabel metal3 s 1821 777 1827 783 3 FreeSans 24 0 0 0 Y[6]
port 8 nsew
flabel metal3 s 1821 737 1827 743 3 FreeSans 24 0 0 0 Y[7]
port 9 nsew
flabel metal2 s 1117 1437 1123 1443 3 FreeSans 24 90 0 0 Y[8]
port 10 nsew
flabel metal2 s 1053 1437 1059 1443 3 FreeSans 24 90 0 0 Y[9]
port 11 nsew
flabel metal2 s 1213 -23 1219 -17 7 FreeSans 24 270 0 0 Y[10]
port 12 nsew
flabel metal2 s 1517 -23 1523 -17 7 FreeSans 24 270 0 0 Y[11]
port 13 nsew
flabel metal2 s 1005 -23 1011 -17 7 FreeSans 24 270 0 0 Y[12]
port 14 nsew
flabel metal2 s 1053 -23 1059 -17 7 FreeSans 24 270 0 0 Y[13]
port 15 nsew
flabel metal2 s 653 -23 659 -17 7 FreeSans 24 270 0 0 Y[14]
port 16 nsew
flabel metal2 s 605 -23 611 -17 7 FreeSans 24 270 0 0 Y[15]
port 17 nsew
flabel metal3 s -19 577 -13 583 7 FreeSans 24 0 0 0 Y[16]
port 18 nsew
flabel metal2 s 381 -23 387 -17 7 FreeSans 24 270 0 0 Y[17]
port 19 nsew
flabel metal3 s -19 657 -13 663 7 FreeSans 24 0 0 0 Y[18]
port 20 nsew
flabel metal3 s -19 697 -13 703 7 FreeSans 24 0 0 0 Y[19]
port 21 nsew
flabel metal3 s -19 1057 -13 1063 7 FreeSans 24 0 0 0 Y[20]
port 22 nsew
flabel metal3 s -19 937 -13 943 7 FreeSans 24 0 0 0 Y[21]
port 23 nsew
flabel metal3 s -19 897 -13 903 7 FreeSans 24 0 0 0 Y[22]
port 24 nsew
flabel metal3 s -19 1097 -13 1103 7 FreeSans 24 0 0 0 Y[23]
port 25 nsew
flabel metal2 s 237 1437 243 1443 3 FreeSans 24 90 0 0 Y[24]
port 26 nsew
flabel metal2 s 189 1437 195 1443 3 FreeSans 24 90 0 0 Y[25]
port 27 nsew
flabel metal2 s 637 1437 643 1443 3 FreeSans 24 90 0 0 Y[26]
port 28 nsew
flabel metal2 s 413 1437 419 1443 3 FreeSans 24 90 0 0 Y[27]
port 29 nsew
flabel metal2 s 925 1437 931 1443 3 FreeSans 24 90 0 0 Y[28]
port 30 nsew
flabel metal2 s 861 1437 867 1443 3 FreeSans 24 90 0 0 Y[29]
port 31 nsew
flabel metal2 s 893 1437 899 1443 3 FreeSans 24 90 0 0 Y[30]
port 32 nsew
flabel metal3 s 1821 697 1827 703 3 FreeSans 24 0 0 0 Y[31]
port 33 nsew
flabel metal2 s 1485 1437 1491 1443 3 FreeSans 24 90 0 0 O[0]
port 34 nsew
flabel metal3 s 1821 1157 1827 1163 3 FreeSans 24 0 0 0 O[1]
port 35 nsew
flabel metal2 s 1469 -23 1475 -17 7 FreeSans 24 270 0 0 O[2]
port 36 nsew
flabel metal3 s 1821 537 1827 543 3 FreeSans 24 0 0 0 O[3]
port 37 nsew
flabel metal2 s 1373 1437 1379 1443 3 FreeSans 24 90 0 0 O[4]
port 38 nsew
flabel metal2 s 1325 1437 1331 1443 3 FreeSans 24 90 0 0 O[5]
port 39 nsew
flabel metal2 s 1405 -23 1411 -17 7 FreeSans 24 270 0 0 O[6]
port 40 nsew
flabel metal2 s 1757 -23 1763 -17 7 FreeSans 24 270 0 0 O[7]
port 41 nsew
flabel metal2 s 941 -23 947 -17 7 FreeSans 24 270 0 0 O[8]
port 42 nsew
flabel metal2 s 1645 -23 1651 -17 7 FreeSans 24 270 0 0 O[9]
port 43 nsew
flabel metal2 s 973 -23 979 -17 7 FreeSans 24 270 0 0 O[10]
port 44 nsew
flabel metal2 s 349 -23 355 -17 7 FreeSans 24 270 0 0 O[11]
port 45 nsew
flabel metal3 s -19 97 -13 103 7 FreeSans 24 0 0 0 O[12]
port 46 nsew
flabel metal2 s 189 -23 195 -17 7 FreeSans 24 270 0 0 O[13]
port 47 nsew
flabel metal2 s 573 -23 579 -17 7 FreeSans 24 270 0 0 O[14]
port 48 nsew
flabel metal3 s 1821 497 1827 503 3 FreeSans 24 0 0 0 O[15]
port 49 nsew
flabel metal3 s -19 137 -13 143 7 FreeSans 24 0 0 0 O[16]
port 50 nsew
flabel metal3 s 1821 1017 1827 1023 3 FreeSans 24 0 0 0 O[17]
port 51 nsew
flabel metal2 s 1581 1437 1587 1443 3 FreeSans 24 90 0 0 O[18]
port 52 nsew
flabel metal3 s -19 1297 -13 1303 7 FreeSans 24 0 0 0 O[19]
port 53 nsew
flabel metal3 s 1821 297 1827 303 3 FreeSans 24 0 0 0 O[20]
port 54 nsew
flabel metal3 s 1821 897 1827 903 3 FreeSans 24 0 0 0 O[21]
port 55 nsew
flabel metal3 s -19 497 -13 503 7 FreeSans 24 0 0 0 O[22]
port 56 nsew
flabel metal3 s -19 537 -13 543 7 FreeSans 24 0 0 0 O[23]
port 57 nsew
flabel metal3 s 1821 817 1827 823 3 FreeSans 24 0 0 0 O[24]
port 58 nsew
flabel metal2 s 1533 1437 1539 1443 3 FreeSans 24 90 0 0 O[25]
port 59 nsew
flabel metal3 s 1821 857 1827 863 3 FreeSans 24 0 0 0 O[26]
port 60 nsew
flabel metal3 s -19 737 -13 743 7 FreeSans 24 0 0 0 O[27]
port 61 nsew
flabel metal2 s 1629 1437 1635 1443 3 FreeSans 24 90 0 0 O[28]
port 62 nsew
flabel metal2 s 1725 1437 1731 1443 3 FreeSans 24 90 0 0 O[29]
port 63 nsew
flabel metal2 s 1421 1437 1427 1443 3 FreeSans 24 90 0 0 O[30]
port 64 nsew
flabel metal2 s 1677 1437 1683 1443 3 FreeSans 24 90 0 0 O[31]
port 65 nsew
<< end >>
