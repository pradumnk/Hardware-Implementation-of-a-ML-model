VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sigmoid_approx
  CLASS BLOCK ;
  FOREIGN sigmoid_approx ;
  ORIGIN 1.900 4.000 ;
  SIZE 184.600 BY 148.300 ;
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 2.800 121.600 3.600 129.000 ;
        RECT 7.600 121.600 8.400 129.800 ;
        RECT 10.800 121.600 11.600 126.200 ;
        RECT 13.000 121.600 13.800 126.200 ;
        RECT 17.200 121.600 18.000 130.200 ;
        RECT 22.000 121.600 22.800 130.200 ;
        RECT 25.800 121.600 26.600 130.200 ;
        RECT 30.000 121.600 30.800 126.200 ;
        RECT 33.200 121.600 34.000 130.200 ;
        RECT 37.400 121.600 38.200 126.200 ;
        RECT 42.200 121.600 43.000 130.200 ;
        RECT 46.000 121.600 46.800 130.200 ;
        RECT 65.200 121.600 66.000 128.200 ;
        RECT 68.400 121.600 69.200 126.200 ;
        RECT 74.800 121.600 75.600 129.000 ;
        RECT 78.000 121.600 78.800 130.200 ;
        RECT 84.400 121.600 85.200 130.200 ;
        RECT 87.600 121.600 88.400 129.000 ;
        RECT 94.000 121.600 94.800 126.200 ;
        RECT 97.200 122.200 98.200 128.800 ;
        RECT 97.400 121.600 98.200 122.200 ;
        RECT 103.400 121.600 104.400 128.800 ;
        RECT 110.000 121.600 110.800 130.200 ;
        RECT 113.200 121.600 114.000 126.200 ;
        RECT 124.400 121.600 125.200 128.200 ;
        RECT 134.000 121.600 134.800 129.000 ;
        RECT 138.800 121.600 139.600 129.000 ;
        RECT 143.600 121.600 144.400 129.000 ;
        RECT 148.400 121.600 149.200 129.000 ;
        RECT 153.200 121.600 154.000 129.000 ;
        RECT 158.000 121.600 158.800 129.000 ;
        RECT 162.800 121.600 163.600 129.000 ;
        RECT 167.600 121.600 168.400 129.000 ;
        RECT 172.400 121.600 173.200 129.000 ;
        RECT 178.800 121.600 179.600 130.200 ;
        RECT 0.400 120.400 180.400 121.600 ;
        RECT 1.200 115.800 2.000 120.400 ;
        RECT 4.400 115.800 5.200 120.400 ;
        RECT 9.200 111.800 10.000 120.400 ;
        RECT 10.800 115.800 11.600 120.400 ;
        RECT 14.600 115.800 15.400 120.400 ;
        RECT 18.800 111.800 19.600 120.400 ;
        RECT 20.400 115.800 21.200 120.400 ;
        RECT 23.600 112.200 24.400 120.400 ;
        RECT 28.400 113.200 29.400 120.400 ;
        RECT 34.600 119.800 35.400 120.400 ;
        RECT 34.600 113.200 35.600 119.800 ;
        RECT 39.600 113.000 40.400 120.400 ;
        RECT 52.400 113.000 53.200 120.400 ;
        RECT 57.200 115.800 58.000 120.400 ;
        RECT 60.400 115.800 61.200 120.400 ;
        RECT 62.600 115.800 63.400 120.400 ;
        RECT 66.800 111.800 67.600 120.400 ;
        RECT 68.400 115.800 69.200 120.400 ;
        RECT 71.600 115.800 72.400 120.400 ;
        RECT 74.800 112.200 75.600 120.400 ;
        RECT 78.000 115.800 78.800 120.400 ;
        RECT 79.600 111.800 80.400 120.400 ;
        RECT 84.400 115.800 85.200 120.400 ;
        RECT 87.600 115.800 88.400 120.400 ;
        RECT 89.200 111.800 90.000 120.400 ;
        RECT 94.000 111.800 94.800 120.400 ;
        RECT 98.200 115.800 99.000 120.400 ;
        RECT 102.200 119.800 103.000 120.400 ;
        RECT 102.000 113.200 103.000 119.800 ;
        RECT 108.200 113.200 109.200 120.400 ;
        RECT 121.200 113.800 122.000 120.400 ;
        RECT 138.800 113.800 139.600 120.400 ;
        RECT 151.600 113.800 152.400 120.400 ;
        RECT 154.800 115.800 155.600 120.400 ;
        RECT 158.000 115.800 158.800 120.400 ;
        RECT 161.200 112.200 162.000 120.400 ;
        RECT 164.400 115.800 165.200 120.400 ;
        RECT 167.600 113.000 168.400 120.400 ;
        RECT 170.800 111.800 171.600 120.400 ;
        RECT 1.200 81.600 2.000 90.200 ;
        RECT 6.000 81.600 6.800 86.200 ;
        RECT 9.200 81.600 10.000 89.800 ;
        RECT 13.600 81.600 14.400 90.200 ;
        RECT 18.800 81.600 19.600 89.800 ;
        RECT 22.000 81.600 22.800 90.200 ;
        RECT 26.200 81.600 27.000 86.200 ;
        RECT 30.000 82.200 31.000 88.800 ;
        RECT 30.200 81.600 31.000 82.200 ;
        RECT 36.200 81.600 37.200 88.800 ;
        RECT 39.600 81.600 40.400 86.200 ;
        RECT 42.800 81.600 43.600 86.200 ;
        RECT 46.000 81.600 46.800 85.800 ;
        RECT 55.600 81.600 56.400 85.800 ;
        RECT 58.800 81.600 59.600 86.200 ;
        RECT 60.400 81.600 61.200 86.200 ;
        RECT 63.600 81.600 64.400 86.200 ;
        RECT 65.200 81.600 66.000 86.200 ;
        RECT 68.400 81.600 69.200 85.800 ;
        RECT 81.200 81.600 82.000 88.200 ;
        RECT 86.000 81.600 86.800 86.200 ;
        RECT 90.800 81.600 91.600 90.200 ;
        RECT 94.000 81.600 94.800 88.200 ;
        RECT 105.800 81.600 106.600 86.200 ;
        RECT 110.000 81.600 110.800 90.200 ;
        RECT 111.600 81.600 112.400 90.200 ;
        RECT 118.000 81.600 118.800 89.000 ;
        RECT 121.200 81.600 122.000 86.200 ;
        RECT 124.400 81.600 125.200 86.200 ;
        RECT 132.400 82.200 133.400 88.800 ;
        RECT 132.600 81.600 133.400 82.200 ;
        RECT 138.600 81.600 139.600 88.800 ;
        RECT 142.600 81.600 143.400 86.200 ;
        RECT 146.800 81.600 147.600 90.200 ;
        RECT 148.400 81.600 149.200 86.200 ;
        RECT 151.600 81.600 152.400 86.200 ;
        RECT 153.200 81.600 154.000 86.200 ;
        RECT 156.400 81.600 157.200 86.200 ;
        RECT 158.000 81.600 158.800 86.200 ;
        RECT 161.200 81.600 162.000 86.200 ;
        RECT 164.400 82.200 165.400 88.800 ;
        RECT 164.600 81.600 165.400 82.200 ;
        RECT 170.600 81.600 171.600 88.800 ;
        RECT 175.600 81.600 176.400 89.000 ;
        RECT 0.400 80.400 180.400 81.600 ;
        RECT 2.800 73.000 3.600 80.400 ;
        RECT 9.200 71.800 10.000 80.400 ;
        RECT 14.000 71.800 14.800 80.400 ;
        RECT 17.200 76.200 18.000 80.400 ;
        RECT 20.400 75.800 21.200 80.400 ;
        RECT 22.000 75.800 22.800 80.400 ;
        RECT 25.200 76.200 26.000 80.400 ;
        RECT 30.000 76.200 30.800 80.400 ;
        RECT 33.200 75.800 34.000 80.400 ;
        RECT 36.400 73.200 37.400 80.400 ;
        RECT 42.600 79.800 43.400 80.400 ;
        RECT 42.600 73.200 43.600 79.800 ;
        RECT 51.400 75.800 52.200 80.400 ;
        RECT 55.600 71.800 56.400 80.400 ;
        RECT 60.400 73.000 61.200 80.400 ;
        RECT 63.600 75.800 64.400 80.400 ;
        RECT 66.800 75.800 67.600 80.400 ;
        RECT 70.000 76.200 70.800 80.400 ;
        RECT 73.200 75.800 74.000 80.400 ;
        RECT 76.400 75.800 77.200 80.400 ;
        RECT 79.600 73.000 80.400 80.400 ;
        RECT 86.000 75.800 86.800 80.400 ;
        RECT 89.200 76.200 90.000 80.400 ;
        RECT 94.000 75.800 94.800 80.400 ;
        RECT 97.200 73.200 98.200 80.400 ;
        RECT 103.400 79.800 104.200 80.400 ;
        RECT 103.400 73.200 104.400 79.800 ;
        RECT 107.400 75.800 108.200 80.400 ;
        RECT 111.600 71.800 112.400 80.400 ;
        RECT 114.800 73.000 115.600 80.400 ;
        RECT 119.600 73.000 120.400 80.400 ;
        RECT 124.400 73.000 125.200 80.400 ;
        RECT 134.000 73.000 134.800 80.400 ;
        RECT 137.200 75.800 138.000 80.400 ;
        RECT 140.400 75.800 141.200 80.400 ;
        RECT 142.600 75.800 143.400 80.400 ;
        RECT 146.800 71.800 147.600 80.400 ;
        RECT 150.200 79.800 151.000 80.400 ;
        RECT 150.000 73.200 151.000 79.800 ;
        RECT 156.200 73.200 157.200 80.400 ;
        RECT 159.600 71.800 160.400 80.400 ;
        RECT 166.000 73.000 166.800 80.400 ;
        RECT 170.800 73.000 171.600 80.400 ;
        RECT 175.600 73.000 176.400 80.400 ;
        RECT 2.800 41.600 3.600 49.000 ;
        RECT 7.600 41.600 8.400 49.000 ;
        RECT 10.800 41.600 11.600 46.200 ;
        RECT 14.000 41.600 14.800 46.200 ;
        RECT 15.600 41.600 16.400 46.200 ;
        RECT 18.800 41.600 19.600 49.800 ;
        RECT 23.600 41.600 24.600 48.800 ;
        RECT 29.800 42.200 30.800 48.800 ;
        RECT 29.800 41.600 30.600 42.200 ;
        RECT 36.400 41.600 37.200 50.200 ;
        RECT 41.200 41.600 42.000 49.000 ;
        RECT 44.400 41.600 45.200 46.200 ;
        RECT 52.400 41.600 53.200 46.200 ;
        RECT 55.600 41.600 56.400 45.800 ;
        RECT 58.800 41.600 59.600 50.200 ;
        RECT 63.000 41.600 63.800 46.200 ;
        RECT 65.200 41.600 66.000 46.200 ;
        RECT 68.400 41.600 69.200 46.200 ;
        RECT 71.600 41.600 72.400 46.200 ;
        RECT 76.400 41.600 77.200 50.200 ;
        RECT 79.600 41.600 80.400 49.000 ;
        RECT 82.800 41.600 83.600 46.200 ;
        RECT 86.000 41.600 86.800 46.200 ;
        RECT 97.200 41.600 98.000 48.200 ;
        RECT 100.400 41.600 101.200 46.200 ;
        RECT 103.600 41.600 104.400 46.200 ;
        RECT 106.800 41.600 107.600 49.800 ;
        RECT 110.000 41.600 110.800 46.200 ;
        RECT 111.600 41.600 112.400 46.200 ;
        RECT 114.800 41.600 115.600 46.200 ;
        RECT 116.400 41.600 117.200 46.200 ;
        RECT 119.600 41.600 120.400 46.200 ;
        RECT 122.800 41.600 123.600 49.000 ;
        RECT 132.400 41.600 133.200 49.000 ;
        RECT 138.800 41.600 139.600 50.200 ;
        RECT 142.000 42.200 143.000 48.800 ;
        RECT 142.200 41.600 143.000 42.200 ;
        RECT 148.200 41.600 149.200 48.800 ;
        RECT 153.200 41.600 154.000 48.200 ;
        RECT 166.000 41.600 166.800 49.000 ;
        RECT 170.800 41.600 171.600 49.000 ;
        RECT 174.000 41.600 174.800 50.200 ;
        RECT 0.400 40.400 180.400 41.600 ;
        RECT 10.800 33.800 11.600 40.400 ;
        RECT 16.200 31.800 17.000 40.400 ;
        RECT 20.400 31.800 21.200 40.400 ;
        RECT 24.600 35.800 25.400 40.400 ;
        RECT 28.400 35.800 29.200 40.400 ;
        RECT 31.600 36.200 32.400 40.400 ;
        RECT 34.800 35.800 35.600 40.400 ;
        RECT 39.600 33.000 40.400 40.400 ;
        RECT 44.600 39.800 45.400 40.400 ;
        RECT 44.400 33.200 45.400 39.800 ;
        RECT 50.600 33.200 51.600 40.400 ;
        RECT 68.400 33.800 69.200 40.400 ;
        RECT 71.600 35.800 72.400 40.400 ;
        RECT 74.800 31.800 75.600 40.400 ;
        RECT 79.000 35.800 79.800 40.400 ;
        RECT 82.800 33.200 83.800 40.400 ;
        RECT 89.000 39.800 89.800 40.400 ;
        RECT 89.000 33.200 90.000 39.800 ;
        RECT 94.000 33.000 94.800 40.400 ;
        RECT 97.200 35.800 98.000 40.400 ;
        RECT 100.400 31.800 101.200 40.400 ;
        RECT 104.600 35.800 105.400 40.400 ;
        RECT 106.800 31.800 107.600 40.400 ;
        RECT 111.000 35.800 111.800 40.400 ;
        RECT 113.200 35.800 114.000 40.400 ;
        RECT 116.400 35.800 117.200 40.400 ;
        RECT 118.000 31.800 118.800 40.400 ;
        RECT 127.600 31.800 128.400 40.400 ;
        RECT 131.800 35.800 132.600 40.400 ;
        RECT 143.600 33.800 144.400 40.400 ;
        RECT 148.600 39.800 149.400 40.400 ;
        RECT 148.400 33.200 149.400 39.800 ;
        RECT 154.600 33.200 155.600 40.400 ;
        RECT 159.600 33.800 160.400 40.400 ;
        RECT 172.400 33.000 173.200 40.400 ;
        RECT 2.800 1.600 3.600 9.000 ;
        RECT 7.600 1.600 8.400 9.000 ;
        RECT 12.400 1.600 13.200 9.800 ;
        RECT 15.600 1.600 16.400 6.200 ;
        RECT 18.800 1.600 19.600 9.000 ;
        RECT 23.600 1.600 24.400 8.200 ;
        RECT 36.400 1.600 37.200 9.000 ;
        RECT 41.200 1.600 42.000 8.200 ;
        RECT 58.800 1.600 59.600 9.000 ;
        RECT 65.200 1.600 66.000 10.200 ;
        RECT 68.400 1.600 69.200 9.800 ;
        RECT 71.600 1.600 72.400 6.200 ;
        RECT 73.200 1.600 74.000 6.200 ;
        RECT 76.400 1.600 77.200 6.200 ;
        RECT 87.600 1.600 88.400 8.200 ;
        RECT 92.400 1.600 93.200 9.000 ;
        RECT 95.600 1.600 96.400 10.200 ;
        RECT 102.000 1.600 103.000 8.800 ;
        RECT 108.200 2.200 109.200 8.800 ;
        RECT 113.200 2.200 114.200 8.800 ;
        RECT 108.200 1.600 109.000 2.200 ;
        RECT 113.400 1.600 114.200 2.200 ;
        RECT 119.400 1.600 120.400 8.800 ;
        RECT 137.200 1.600 138.000 8.200 ;
        RECT 142.000 1.600 142.800 9.000 ;
        RECT 146.800 1.600 147.600 9.000 ;
        RECT 159.600 1.600 160.400 8.200 ;
        RECT 164.400 1.600 165.200 9.000 ;
        RECT 169.200 1.600 170.000 9.800 ;
        RECT 172.400 1.600 173.200 6.200 ;
        RECT 175.600 1.600 176.400 9.000 ;
        RECT 0.400 0.400 180.400 1.600 ;
      LAYER via1 ;
        RECT 49.400 120.600 50.200 121.400 ;
        RECT 50.800 120.600 51.600 121.400 ;
        RECT 52.200 120.600 53.000 121.400 ;
        RECT 49.400 80.600 50.200 81.400 ;
        RECT 50.800 80.600 51.600 81.400 ;
        RECT 52.200 80.600 53.000 81.400 ;
        RECT 49.400 40.600 50.200 41.400 ;
        RECT 50.800 40.600 51.600 41.400 ;
        RECT 52.200 40.600 53.000 41.400 ;
        RECT 49.400 0.600 50.200 1.400 ;
        RECT 50.800 0.600 51.600 1.400 ;
        RECT 52.200 0.600 53.000 1.400 ;
      LAYER metal2 ;
        RECT 48.800 120.600 53.600 121.400 ;
        RECT 48.800 80.600 53.600 81.400 ;
        RECT 48.800 40.600 53.600 41.400 ;
        RECT 48.800 0.600 53.600 1.400 ;
      LAYER via2 ;
        RECT 49.400 120.600 50.200 121.400 ;
        RECT 50.800 120.600 51.600 121.400 ;
        RECT 52.200 120.600 53.000 121.400 ;
        RECT 49.400 80.600 50.200 81.400 ;
        RECT 50.800 80.600 51.600 81.400 ;
        RECT 52.200 80.600 53.000 81.400 ;
        RECT 49.400 40.600 50.200 41.400 ;
        RECT 50.800 40.600 51.600 41.400 ;
        RECT 52.200 40.600 53.000 41.400 ;
        RECT 49.400 0.600 50.200 1.400 ;
        RECT 50.800 0.600 51.600 1.400 ;
        RECT 52.200 0.600 53.000 1.400 ;
      LAYER metal3 ;
        RECT 48.800 120.400 53.600 121.600 ;
        RECT 48.800 80.400 53.600 81.600 ;
        RECT 48.800 40.400 53.600 41.600 ;
        RECT 48.800 0.400 53.600 1.600 ;
      LAYER via3 ;
        RECT 49.200 120.600 50.000 121.400 ;
        RECT 50.800 120.600 51.600 121.400 ;
        RECT 52.400 120.600 53.200 121.400 ;
        RECT 49.200 80.600 50.000 81.400 ;
        RECT 50.800 80.600 51.600 81.400 ;
        RECT 52.400 80.600 53.200 81.400 ;
        RECT 49.200 40.600 50.000 41.400 ;
        RECT 50.800 40.600 51.600 41.400 ;
        RECT 52.400 40.600 53.200 41.400 ;
        RECT 49.200 0.600 50.000 1.400 ;
        RECT 50.800 0.600 51.600 1.400 ;
        RECT 52.400 0.600 53.200 1.400 ;
      LAYER metal4 ;
        RECT 48.800 -4.000 53.600 144.000 ;
    END
  END vdd
  PIN gnd
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.400 140.400 180.400 141.600 ;
        RECT 2.800 135.800 3.600 140.400 ;
        RECT 8.200 136.000 9.000 140.400 ;
        RECT 15.600 136.600 16.400 140.400 ;
        RECT 18.800 137.800 19.600 140.400 ;
        RECT 22.000 137.800 22.800 140.400 ;
        RECT 25.200 136.200 26.000 140.400 ;
        RECT 28.400 137.800 29.200 140.400 ;
        RECT 30.000 137.800 30.800 140.400 ;
        RECT 34.800 136.600 35.600 140.400 ;
        RECT 39.600 137.800 40.400 140.400 ;
        RECT 42.800 136.200 43.600 140.400 ;
        RECT 46.000 137.800 46.800 140.400 ;
        RECT 49.200 137.800 50.000 140.400 ;
        RECT 62.000 138.200 62.800 140.400 ;
        RECT 65.200 137.800 66.000 140.400 ;
        RECT 68.400 137.800 69.200 140.400 ;
        RECT 71.600 137.800 72.400 140.400 ;
        RECT 75.800 135.800 76.600 140.400 ;
        RECT 79.600 136.600 80.400 140.400 ;
        RECT 86.600 135.800 87.400 140.400 ;
        RECT 90.800 137.800 91.600 140.400 ;
        RECT 94.000 137.800 94.800 140.400 ;
        RECT 97.400 139.800 98.200 140.400 ;
        RECT 97.200 136.400 98.200 139.800 ;
        RECT 103.400 136.400 104.400 140.400 ;
        RECT 106.800 137.800 107.600 140.400 ;
        RECT 110.000 137.800 110.800 140.400 ;
        RECT 113.200 137.800 114.000 140.400 ;
        RECT 121.200 138.200 122.000 140.400 ;
        RECT 124.400 137.800 125.200 140.400 ;
        RECT 134.000 135.800 134.800 140.400 ;
        RECT 138.800 135.800 139.600 140.400 ;
        RECT 143.600 135.800 144.400 140.400 ;
        RECT 148.400 135.800 149.200 140.400 ;
        RECT 153.200 135.800 154.000 140.400 ;
        RECT 158.000 135.800 158.800 140.400 ;
        RECT 162.800 135.800 163.600 140.400 ;
        RECT 167.600 135.800 168.400 140.400 ;
        RECT 172.400 135.800 173.200 140.400 ;
        RECT 175.600 137.800 176.400 140.400 ;
        RECT 178.800 137.800 179.600 140.400 ;
        RECT 4.400 131.600 5.200 133.200 ;
        RECT 142.000 131.600 142.800 133.200 ;
        RECT 151.600 131.600 152.400 133.200 ;
        RECT 156.400 131.600 157.200 133.200 ;
        RECT 161.200 131.600 162.000 133.200 ;
        RECT 166.000 131.600 166.800 133.200 ;
        RECT 170.800 131.600 171.600 133.200 ;
        RECT 1.200 101.600 2.000 106.200 ;
        RECT 6.000 101.600 6.800 104.200 ;
        RECT 9.200 101.600 10.000 104.200 ;
        RECT 10.800 101.600 11.600 104.200 ;
        RECT 17.200 101.600 18.000 105.400 ;
        RECT 23.000 101.600 23.800 106.000 ;
        RECT 28.400 101.600 29.400 105.600 ;
        RECT 34.600 102.200 35.600 105.600 ;
        RECT 34.600 101.600 35.400 102.200 ;
        RECT 38.400 101.600 39.200 106.200 ;
        RECT 44.400 101.600 45.200 106.200 ;
        RECT 51.400 101.600 52.200 106.200 ;
        RECT 55.600 101.600 56.400 104.200 ;
        RECT 57.200 101.600 58.000 106.200 ;
        RECT 65.200 101.600 66.000 105.400 ;
        RECT 71.600 101.600 72.400 106.200 ;
        RECT 75.400 101.600 76.200 106.000 ;
        RECT 79.600 101.600 80.400 104.200 ;
        RECT 82.800 101.600 83.600 104.200 ;
        RECT 87.600 101.600 88.400 106.200 ;
        RECT 89.200 101.600 90.000 104.200 ;
        RECT 92.400 101.600 93.200 104.200 ;
        RECT 95.600 101.600 96.400 105.400 ;
        RECT 102.000 102.200 103.000 105.600 ;
        RECT 102.200 101.600 103.000 102.200 ;
        RECT 108.200 101.600 109.200 105.600 ;
        RECT 118.000 101.600 118.800 103.800 ;
        RECT 121.200 101.600 122.000 104.200 ;
        RECT 135.600 101.600 136.400 103.800 ;
        RECT 138.800 101.600 139.600 104.200 ;
        RECT 148.400 101.600 149.200 103.800 ;
        RECT 151.600 101.600 152.400 104.200 ;
        RECT 158.000 101.600 158.800 106.200 ;
        RECT 161.800 101.600 162.600 106.000 ;
        RECT 167.600 101.600 168.400 106.200 ;
        RECT 170.800 101.600 171.600 104.200 ;
        RECT 174.000 101.600 174.800 104.200 ;
        RECT 0.400 100.400 180.400 101.600 ;
        RECT 1.200 97.800 2.000 100.400 ;
        RECT 4.400 97.800 5.200 100.400 ;
        RECT 8.600 96.000 9.400 100.400 ;
        RECT 13.600 95.000 14.400 100.400 ;
        RECT 18.800 95.400 19.600 100.400 ;
        RECT 23.600 96.600 24.400 100.400 ;
        RECT 30.200 99.800 31.000 100.400 ;
        RECT 30.000 96.400 31.000 99.800 ;
        RECT 36.200 96.400 37.200 100.400 ;
        RECT 39.600 97.800 40.400 100.400 ;
        RECT 42.800 93.800 43.600 100.400 ;
        RECT 58.800 93.800 59.600 100.400 ;
        RECT 60.400 95.800 61.200 100.400 ;
        RECT 65.200 93.800 66.000 100.400 ;
        RECT 78.000 98.200 78.800 100.400 ;
        RECT 81.200 97.800 82.000 100.400 ;
        RECT 86.000 97.800 86.800 100.400 ;
        RECT 87.600 97.800 88.400 100.400 ;
        RECT 90.800 97.800 91.600 100.400 ;
        RECT 94.000 97.800 94.800 100.400 ;
        RECT 97.200 98.200 98.000 100.400 ;
        RECT 108.400 96.600 109.200 100.400 ;
        RECT 111.600 97.800 112.400 100.400 ;
        RECT 114.800 97.800 115.600 100.400 ;
        RECT 118.000 95.800 118.800 100.400 ;
        RECT 121.200 95.800 122.000 100.400 ;
        RECT 132.600 99.800 133.400 100.400 ;
        RECT 132.400 96.400 133.400 99.800 ;
        RECT 138.600 96.400 139.600 100.400 ;
        RECT 145.200 96.600 146.000 100.400 ;
        RECT 151.600 95.800 152.400 100.400 ;
        RECT 153.200 95.800 154.000 100.400 ;
        RECT 158.000 95.800 158.800 100.400 ;
        RECT 164.600 99.800 165.400 100.400 ;
        RECT 164.400 96.400 165.400 99.800 ;
        RECT 170.600 96.400 171.600 100.400 ;
        RECT 175.600 95.800 176.400 100.400 ;
        RECT 174.000 91.600 174.800 93.200 ;
        RECT 4.400 68.800 5.200 70.400 ;
        RECT 167.600 70.300 168.400 70.400 ;
        RECT 169.200 70.300 170.000 70.400 ;
        RECT 167.600 69.700 170.000 70.300 ;
        RECT 167.600 68.800 168.400 69.700 ;
        RECT 169.200 68.800 170.000 69.700 ;
        RECT 174.000 68.800 174.800 70.400 ;
        RECT 2.800 61.600 3.600 66.200 ;
        RECT 6.000 61.600 6.800 64.200 ;
        RECT 9.200 61.600 10.000 64.200 ;
        RECT 10.800 61.600 11.600 64.200 ;
        RECT 14.000 61.600 14.800 64.200 ;
        RECT 20.400 61.600 21.200 68.200 ;
        RECT 22.000 61.600 22.800 68.200 ;
        RECT 33.200 61.600 34.000 68.200 ;
        RECT 36.400 61.600 37.400 65.600 ;
        RECT 42.600 62.200 43.600 65.600 ;
        RECT 42.600 61.600 43.400 62.200 ;
        RECT 54.000 61.600 54.800 65.400 ;
        RECT 57.200 61.600 58.000 64.200 ;
        RECT 61.400 61.600 62.200 66.200 ;
        RECT 63.600 61.600 64.400 64.200 ;
        RECT 66.800 61.600 67.600 68.200 ;
        RECT 76.400 61.600 77.200 66.200 ;
        RECT 78.400 61.600 79.200 66.200 ;
        RECT 84.400 61.600 85.200 66.200 ;
        RECT 86.000 61.600 86.800 68.200 ;
        RECT 94.000 61.600 94.800 64.200 ;
        RECT 97.200 61.600 98.200 65.600 ;
        RECT 103.400 62.200 104.400 65.600 ;
        RECT 103.400 61.600 104.200 62.200 ;
        RECT 110.000 61.600 110.800 65.400 ;
        RECT 114.800 61.600 115.600 66.200 ;
        RECT 119.600 61.600 120.400 66.200 ;
        RECT 124.400 61.600 125.200 66.200 ;
        RECT 134.000 61.600 134.800 66.200 ;
        RECT 137.200 61.600 138.000 66.200 ;
        RECT 145.200 61.600 146.000 65.400 ;
        RECT 150.000 62.200 151.000 65.600 ;
        RECT 150.200 61.600 151.000 62.200 ;
        RECT 156.200 61.600 157.200 65.600 ;
        RECT 159.600 61.600 160.400 64.200 ;
        RECT 162.800 61.600 163.600 64.200 ;
        RECT 166.000 61.600 166.800 66.200 ;
        RECT 170.800 61.600 171.600 66.200 ;
        RECT 175.600 61.600 176.400 66.200 ;
        RECT 0.400 60.400 180.400 61.600 ;
        RECT 2.800 55.800 3.600 60.400 ;
        RECT 7.600 55.800 8.400 60.400 ;
        RECT 14.000 55.800 14.800 60.400 ;
        RECT 18.200 56.000 19.000 60.400 ;
        RECT 23.600 56.400 24.600 60.400 ;
        RECT 29.800 59.800 30.600 60.400 ;
        RECT 29.800 56.400 30.800 59.800 ;
        RECT 33.200 57.800 34.000 60.400 ;
        RECT 36.400 57.800 37.200 60.400 ;
        RECT 38.000 57.800 38.800 60.400 ;
        RECT 42.200 55.800 43.000 60.400 ;
        RECT 44.400 57.800 45.200 60.400 ;
        RECT 52.400 53.800 53.200 60.400 ;
        RECT 60.400 56.600 61.200 60.400 ;
        RECT 65.200 55.800 66.000 60.400 ;
        RECT 71.600 57.800 72.400 60.400 ;
        RECT 73.200 57.800 74.000 60.400 ;
        RECT 76.400 57.800 77.200 60.400 ;
        RECT 79.600 55.800 80.400 60.400 ;
        RECT 86.000 55.800 86.800 60.400 ;
        RECT 94.000 58.200 94.800 60.400 ;
        RECT 97.200 57.800 98.000 60.400 ;
        RECT 103.600 55.800 104.400 60.400 ;
        RECT 107.400 56.000 108.200 60.400 ;
        RECT 114.800 55.800 115.600 60.400 ;
        RECT 119.600 55.800 120.400 60.400 ;
        RECT 122.800 55.800 123.600 60.400 ;
        RECT 132.400 55.800 133.200 60.400 ;
        RECT 135.600 57.800 136.400 60.400 ;
        RECT 138.800 57.800 139.600 60.400 ;
        RECT 142.200 59.800 143.000 60.400 ;
        RECT 142.000 56.400 143.000 59.800 ;
        RECT 148.200 56.400 149.200 60.400 ;
        RECT 153.200 57.800 154.000 60.400 ;
        RECT 156.400 58.200 157.200 60.400 ;
        RECT 166.000 55.800 166.800 60.400 ;
        RECT 170.800 55.800 171.600 60.400 ;
        RECT 174.000 57.800 174.800 60.400 ;
        RECT 177.200 57.800 178.000 60.400 ;
        RECT 4.400 51.600 5.200 53.200 ;
        RECT 9.200 51.600 10.000 53.200 ;
        RECT 170.800 28.800 171.600 30.400 ;
        RECT 7.600 21.600 8.400 23.800 ;
        RECT 10.800 21.600 11.600 24.200 ;
        RECT 15.600 21.600 16.400 25.800 ;
        RECT 18.800 21.600 19.600 24.200 ;
        RECT 22.000 21.600 22.800 25.400 ;
        RECT 28.400 21.600 29.200 24.200 ;
        RECT 34.800 21.600 35.600 28.200 ;
        RECT 36.400 21.600 37.200 24.200 ;
        RECT 40.600 21.600 41.400 26.200 ;
        RECT 44.400 22.200 45.400 25.600 ;
        RECT 44.600 21.600 45.400 22.200 ;
        RECT 50.600 21.600 51.600 25.600 ;
        RECT 65.200 21.600 66.000 23.800 ;
        RECT 68.400 21.600 69.200 24.200 ;
        RECT 71.600 21.600 72.400 24.200 ;
        RECT 76.400 21.600 77.200 25.400 ;
        RECT 82.800 21.600 83.800 25.600 ;
        RECT 89.000 22.200 90.000 25.600 ;
        RECT 89.000 21.600 89.800 22.200 ;
        RECT 94.000 21.600 94.800 26.200 ;
        RECT 97.200 21.600 98.000 24.200 ;
        RECT 102.000 21.600 102.800 25.400 ;
        RECT 108.400 21.600 109.200 25.400 ;
        RECT 113.200 21.600 114.000 26.200 ;
        RECT 118.000 21.600 118.800 24.200 ;
        RECT 121.200 21.600 122.000 24.200 ;
        RECT 129.200 21.600 130.000 25.400 ;
        RECT 140.400 21.600 141.200 23.800 ;
        RECT 143.600 21.600 144.400 24.200 ;
        RECT 148.400 22.200 149.400 25.600 ;
        RECT 148.600 21.600 149.400 22.200 ;
        RECT 154.600 21.600 155.600 25.600 ;
        RECT 159.600 21.600 160.400 24.200 ;
        RECT 162.800 21.600 163.600 23.800 ;
        RECT 172.400 21.600 173.200 26.200 ;
        RECT 0.400 20.400 180.400 21.600 ;
        RECT 2.800 15.800 3.600 20.400 ;
        RECT 7.600 15.800 8.400 20.400 ;
        RECT 13.000 16.000 13.800 20.400 ;
        RECT 18.800 15.800 19.600 20.400 ;
        RECT 23.600 17.800 24.400 20.400 ;
        RECT 26.800 18.200 27.600 20.400 ;
        RECT 36.400 15.800 37.200 20.400 ;
        RECT 41.200 17.800 42.000 20.400 ;
        RECT 44.400 18.200 45.200 20.400 ;
        RECT 58.800 15.800 59.600 20.400 ;
        RECT 62.000 17.800 62.800 20.400 ;
        RECT 65.200 17.800 66.000 20.400 ;
        RECT 69.000 16.000 69.800 20.400 ;
        RECT 76.400 15.800 77.200 20.400 ;
        RECT 84.400 18.200 85.200 20.400 ;
        RECT 87.600 17.800 88.400 20.400 ;
        RECT 92.400 15.800 93.200 20.400 ;
        RECT 95.600 17.800 96.400 20.400 ;
        RECT 98.800 17.800 99.600 20.400 ;
        RECT 102.000 16.400 103.000 20.400 ;
        RECT 108.200 19.800 109.000 20.400 ;
        RECT 113.400 19.800 114.200 20.400 ;
        RECT 108.200 16.400 109.200 19.800 ;
        RECT 113.200 16.400 114.200 19.800 ;
        RECT 119.400 16.400 120.400 20.400 ;
        RECT 134.000 18.200 134.800 20.400 ;
        RECT 137.200 17.800 138.000 20.400 ;
        RECT 142.000 15.800 142.800 20.400 ;
        RECT 146.800 15.800 147.600 20.400 ;
        RECT 156.400 18.200 157.200 20.400 ;
        RECT 159.600 17.800 160.400 20.400 ;
        RECT 164.400 15.800 165.200 20.400 ;
        RECT 169.800 16.000 170.600 20.400 ;
        RECT 175.600 15.800 176.400 20.400 ;
      LAYER via1 ;
        RECT 124.600 140.600 125.400 141.400 ;
        RECT 126.000 140.600 126.800 141.400 ;
        RECT 127.400 140.600 128.200 141.400 ;
        RECT 124.600 100.600 125.400 101.400 ;
        RECT 126.000 100.600 126.800 101.400 ;
        RECT 127.400 100.600 128.200 101.400 ;
        RECT 4.400 69.600 5.200 70.400 ;
        RECT 167.600 69.600 168.400 70.400 ;
        RECT 174.000 69.600 174.800 70.400 ;
        RECT 2.800 65.400 3.600 66.200 ;
        RECT 166.000 65.400 166.800 66.200 ;
        RECT 124.600 60.600 125.400 61.400 ;
        RECT 126.000 60.600 126.800 61.400 ;
        RECT 127.400 60.600 128.200 61.400 ;
        RECT 174.000 59.600 174.800 60.400 ;
        RECT 170.800 29.600 171.600 30.400 ;
        RECT 172.400 25.400 173.200 26.200 ;
        RECT 124.600 20.600 125.400 21.400 ;
        RECT 126.000 20.600 126.800 21.400 ;
        RECT 127.400 20.600 128.200 21.400 ;
      LAYER metal2 ;
        RECT 124.000 140.600 128.800 141.400 ;
        RECT 2.800 136.300 3.600 136.600 ;
        RECT 143.600 136.300 144.400 136.600 ;
        RECT 153.200 136.300 154.000 136.600 ;
        RECT 158.000 136.300 158.800 136.600 ;
        RECT 162.800 136.300 163.600 136.600 ;
        RECT 167.600 136.300 168.400 136.600 ;
        RECT 172.400 136.300 173.200 136.600 ;
        RECT 2.800 135.800 5.100 136.300 ;
        RECT 2.900 135.700 5.100 135.800 ;
        RECT 4.500 132.400 5.100 135.700 ;
        RECT 142.100 135.800 144.400 136.300 ;
        RECT 151.700 135.800 154.000 136.300 ;
        RECT 156.500 135.800 158.800 136.300 ;
        RECT 161.300 135.800 163.600 136.300 ;
        RECT 166.100 135.800 168.400 136.300 ;
        RECT 170.900 135.800 173.200 136.300 ;
        RECT 142.100 135.700 144.300 135.800 ;
        RECT 151.700 135.700 153.900 135.800 ;
        RECT 156.500 135.700 158.700 135.800 ;
        RECT 161.300 135.700 163.500 135.800 ;
        RECT 166.100 135.700 168.300 135.800 ;
        RECT 170.900 135.700 173.100 135.800 ;
        RECT 142.100 132.400 142.700 135.700 ;
        RECT 151.700 132.400 152.300 135.700 ;
        RECT 156.500 132.400 157.100 135.700 ;
        RECT 161.300 132.400 161.900 135.700 ;
        RECT 166.100 132.400 166.700 135.700 ;
        RECT 170.900 132.400 171.500 135.700 ;
        RECT 4.400 131.600 5.200 132.400 ;
        RECT 142.000 131.600 142.800 132.400 ;
        RECT 151.600 131.600 152.400 132.400 ;
        RECT 156.400 131.600 157.200 132.400 ;
        RECT 161.200 131.600 162.000 132.400 ;
        RECT 166.000 131.600 166.800 132.400 ;
        RECT 170.800 131.600 171.600 132.400 ;
        RECT 174.000 101.600 174.800 102.400 ;
        RECT 124.000 100.600 128.800 101.400 ;
        RECT 174.100 92.400 174.700 101.600 ;
        RECT 174.000 91.600 174.800 92.400 ;
        RECT 4.400 69.600 5.200 70.400 ;
        RECT 167.600 69.600 168.400 70.400 ;
        RECT 174.000 69.600 174.800 70.400 ;
        RECT 4.500 66.300 5.100 69.600 ;
        RECT 167.700 66.300 168.300 69.600 ;
        RECT 2.900 66.200 5.100 66.300 ;
        RECT 166.100 66.200 168.300 66.300 ;
        RECT 2.800 65.700 5.100 66.200 ;
        RECT 166.000 65.700 168.300 66.200 ;
        RECT 2.800 65.400 3.600 65.700 ;
        RECT 166.000 65.400 166.800 65.700 ;
        RECT 9.200 61.600 10.000 62.400 ;
        RECT 2.800 56.300 3.600 56.600 ;
        RECT 2.800 55.800 5.100 56.300 ;
        RECT 2.900 55.700 5.100 55.800 ;
        RECT 4.500 52.400 5.100 55.700 ;
        RECT 9.300 52.400 9.900 61.600 ;
        RECT 124.000 60.600 128.800 61.400 ;
        RECT 174.100 60.400 174.700 69.600 ;
        RECT 174.000 59.600 174.800 60.400 ;
        RECT 4.400 51.600 5.200 52.400 ;
        RECT 9.200 51.600 10.000 52.400 ;
        RECT 170.800 29.600 171.600 30.400 ;
        RECT 170.900 26.300 171.500 29.600 ;
        RECT 170.900 26.200 173.100 26.300 ;
        RECT 170.900 25.700 173.200 26.200 ;
        RECT 172.400 25.400 173.200 25.700 ;
        RECT 124.000 20.600 128.800 21.400 ;
      LAYER via2 ;
        RECT 124.600 140.600 125.400 141.400 ;
        RECT 126.000 140.600 126.800 141.400 ;
        RECT 127.400 140.600 128.200 141.400 ;
        RECT 124.600 100.600 125.400 101.400 ;
        RECT 126.000 100.600 126.800 101.400 ;
        RECT 127.400 100.600 128.200 101.400 ;
        RECT 124.600 60.600 125.400 61.400 ;
        RECT 126.000 60.600 126.800 61.400 ;
        RECT 127.400 60.600 128.200 61.400 ;
        RECT 124.600 20.600 125.400 21.400 ;
        RECT 126.000 20.600 126.800 21.400 ;
        RECT 127.400 20.600 128.200 21.400 ;
      LAYER metal3 ;
        RECT 124.000 140.400 128.800 141.600 ;
        RECT 124.000 100.400 128.800 101.600 ;
        RECT 124.000 60.400 128.800 61.600 ;
        RECT 124.000 20.400 128.800 21.600 ;
      LAYER via3 ;
        RECT 124.400 140.600 125.200 141.400 ;
        RECT 126.000 140.600 126.800 141.400 ;
        RECT 127.600 140.600 128.400 141.400 ;
        RECT 124.400 100.600 125.200 101.400 ;
        RECT 126.000 100.600 126.800 101.400 ;
        RECT 127.600 100.600 128.400 101.400 ;
        RECT 124.400 60.600 125.200 61.400 ;
        RECT 126.000 60.600 126.800 61.400 ;
        RECT 127.600 60.600 128.400 61.400 ;
        RECT 124.400 20.600 125.200 21.400 ;
        RECT 126.000 20.600 126.800 21.400 ;
        RECT 127.600 20.600 128.400 21.400 ;
      LAYER metal4 ;
        RECT 124.000 -4.000 128.800 144.000 ;
    END
  END gnd
  PIN Y[0]
    PORT
      LAYER metal1 ;
        RECT 170.800 104.800 171.600 106.400 ;
      LAYER via1 ;
        RECT 170.800 105.600 171.600 106.400 ;
      LAYER metal2 ;
        RECT 170.800 105.600 171.600 106.400 ;
      LAYER metal3 ;
        RECT 178.900 107.700 182.700 108.300 ;
        RECT 170.800 106.300 171.600 106.400 ;
        RECT 178.900 106.300 179.500 107.700 ;
        RECT 170.800 105.700 179.500 106.300 ;
        RECT 170.800 105.600 171.600 105.700 ;
    END
  END Y[0]
  PIN Y[1]
    PORT
      LAYER metal1 ;
        RECT 178.800 135.600 179.600 137.200 ;
      LAYER metal2 ;
        RECT 178.900 143.700 181.100 144.300 ;
        RECT 178.900 136.400 179.500 143.700 ;
        RECT 178.800 135.600 179.600 136.400 ;
    END
  END Y[1]
  PIN Y[2]
    PORT
      LAYER metal1 ;
        RECT 175.600 130.800 176.400 132.400 ;
      LAYER via1 ;
        RECT 175.600 131.600 176.400 132.400 ;
      LAYER metal2 ;
        RECT 175.700 143.700 177.900 144.300 ;
        RECT 175.700 132.400 176.300 143.700 ;
        RECT 175.600 131.600 176.400 132.400 ;
    END
  END Y[2]
  PIN Y[3]
    PORT
      LAYER metal1 ;
        RECT 174.000 110.300 174.800 111.200 ;
        RECT 178.800 110.300 179.600 110.400 ;
        RECT 174.000 109.700 179.600 110.300 ;
        RECT 174.000 109.600 174.800 109.700 ;
        RECT 178.800 109.600 179.600 109.700 ;
      LAYER metal2 ;
        RECT 178.800 111.600 179.600 112.400 ;
        RECT 178.900 110.400 179.500 111.600 ;
        RECT 178.800 109.600 179.600 110.400 ;
      LAYER metal3 ;
        RECT 178.800 112.300 179.600 112.400 ;
        RECT 178.800 111.700 182.700 112.300 ;
        RECT 178.800 111.600 179.600 111.700 ;
    END
  END Y[3]
  PIN Y[4]
    PORT
      LAYER metal1 ;
        RECT 146.000 94.400 146.800 94.800 ;
        RECT 139.600 93.600 141.200 94.400 ;
        RECT 146.000 93.800 147.600 94.400 ;
        RECT 146.800 93.600 147.600 93.800 ;
        RECT 177.200 52.300 178.000 52.400 ;
        RECT 178.800 52.300 179.600 52.400 ;
        RECT 177.200 51.700 179.600 52.300 ;
        RECT 177.200 50.800 178.000 51.700 ;
        RECT 178.800 51.600 179.600 51.700 ;
      LAYER via1 ;
        RECT 140.400 93.600 141.200 94.400 ;
      LAYER metal2 ;
        RECT 178.800 95.600 179.600 96.400 ;
        RECT 140.400 93.600 141.200 94.400 ;
        RECT 146.800 93.600 147.600 94.400 ;
        RECT 140.500 86.400 141.100 93.600 ;
        RECT 146.900 86.400 147.500 93.600 ;
        RECT 178.900 86.400 179.500 95.600 ;
        RECT 140.400 85.600 141.200 86.400 ;
        RECT 146.800 85.600 147.600 86.400 ;
        RECT 178.800 85.600 179.600 86.400 ;
        RECT 178.900 52.400 179.500 85.600 ;
        RECT 178.800 51.600 179.600 52.400 ;
      LAYER metal3 ;
        RECT 180.500 97.700 182.700 98.300 ;
        RECT 178.800 96.300 179.600 96.400 ;
        RECT 180.500 96.300 181.100 97.700 ;
        RECT 178.800 95.700 181.100 96.300 ;
        RECT 178.800 95.600 179.600 95.700 ;
        RECT 140.400 86.300 141.200 86.400 ;
        RECT 146.800 86.300 147.600 86.400 ;
        RECT 178.800 86.300 179.600 86.400 ;
        RECT 140.400 85.700 179.600 86.300 ;
        RECT 140.400 85.600 141.200 85.700 ;
        RECT 146.800 85.600 147.600 85.700 ;
        RECT 178.800 85.600 179.600 85.700 ;
    END
  END Y[4]
  PIN Y[5]
    PORT
      LAYER metal1 ;
        RECT 171.600 93.600 173.200 94.400 ;
        RECT 174.000 55.600 174.800 57.200 ;
      LAYER via1 ;
        RECT 172.400 93.600 173.200 94.400 ;
      LAYER metal2 ;
        RECT 172.400 93.600 173.200 94.400 ;
        RECT 174.000 57.600 174.800 58.400 ;
        RECT 174.100 56.400 174.700 57.600 ;
        RECT 174.000 55.600 174.800 56.400 ;
      LAYER metal3 ;
        RECT 172.400 94.300 173.200 94.400 ;
        RECT 174.000 94.300 174.800 94.400 ;
        RECT 172.400 93.700 182.700 94.300 ;
        RECT 172.400 93.600 173.200 93.700 ;
        RECT 174.000 93.600 174.800 93.700 ;
        RECT 174.000 57.600 174.800 58.400 ;
      LAYER metal4 ;
        RECT 173.800 57.400 175.000 94.600 ;
    END
  END Y[5]
  PIN Y[6]
    PORT
      LAYER metal1 ;
        RECT 146.800 68.200 147.600 68.400 ;
        RECT 146.000 67.600 147.600 68.200 ;
        RECT 146.000 67.200 146.800 67.600 ;
        RECT 159.600 64.800 160.400 66.400 ;
        RECT 149.200 53.600 150.800 54.400 ;
      LAYER via1 ;
        RECT 146.800 67.600 147.600 68.400 ;
        RECT 159.600 65.600 160.400 66.400 ;
        RECT 150.000 53.600 150.800 54.400 ;
      LAYER metal2 ;
        RECT 159.600 77.600 160.400 78.400 ;
        RECT 146.800 67.600 147.600 68.400 ;
        RECT 146.900 66.400 147.500 67.600 ;
        RECT 159.700 66.400 160.300 77.600 ;
        RECT 146.800 65.600 147.600 66.400 ;
        RECT 159.600 65.600 160.400 66.400 ;
        RECT 146.900 58.400 147.500 65.600 ;
        RECT 146.800 57.600 147.600 58.400 ;
        RECT 150.000 57.600 150.800 58.400 ;
        RECT 150.100 54.400 150.700 57.600 ;
        RECT 150.000 53.600 150.800 54.400 ;
      LAYER metal3 ;
        RECT 159.600 78.300 160.400 78.400 ;
        RECT 159.600 77.700 182.700 78.300 ;
        RECT 159.600 77.600 160.400 77.700 ;
        RECT 146.800 66.300 147.600 66.400 ;
        RECT 159.600 66.300 160.400 66.400 ;
        RECT 146.800 65.700 160.400 66.300 ;
        RECT 146.800 65.600 147.600 65.700 ;
        RECT 159.600 65.600 160.400 65.700 ;
        RECT 146.800 58.300 147.600 58.400 ;
        RECT 150.000 58.300 150.800 58.400 ;
        RECT 146.800 57.700 150.800 58.300 ;
        RECT 146.800 57.600 147.600 57.700 ;
        RECT 150.000 57.600 150.800 57.700 ;
    END
  END Y[6]
  PIN Y[7]
    PORT
      LAYER metal1 ;
        RECT 162.800 69.600 163.600 71.200 ;
        RECT 157.200 67.600 158.800 68.400 ;
      LAYER via1 ;
        RECT 158.000 67.600 158.800 68.400 ;
      LAYER metal2 ;
        RECT 158.000 73.600 158.800 74.400 ;
        RECT 162.800 73.600 163.600 74.400 ;
        RECT 158.100 68.400 158.700 73.600 ;
        RECT 162.900 70.400 163.500 73.600 ;
        RECT 162.800 69.600 163.600 70.400 ;
        RECT 158.000 67.600 158.800 68.400 ;
      LAYER metal3 ;
        RECT 158.000 74.300 158.800 74.400 ;
        RECT 162.800 74.300 163.600 74.400 ;
        RECT 158.000 73.700 182.700 74.300 ;
        RECT 158.000 73.600 158.800 73.700 ;
        RECT 162.800 73.600 163.600 73.700 ;
    END
  END Y[7]
  PIN Y[8]
    PORT
      LAYER metal1 ;
        RECT 110.000 135.600 110.800 137.200 ;
        RECT 113.200 135.600 114.000 137.200 ;
      LAYER metal2 ;
        RECT 110.100 143.700 112.300 144.300 ;
        RECT 110.100 136.400 110.700 143.700 ;
        RECT 110.000 135.600 110.800 136.400 ;
        RECT 113.200 135.600 114.000 136.400 ;
      LAYER metal3 ;
        RECT 110.000 136.300 110.800 136.400 ;
        RECT 113.200 136.300 114.000 136.400 ;
        RECT 110.000 135.700 114.000 136.300 ;
        RECT 110.000 135.600 110.800 135.700 ;
        RECT 113.200 135.600 114.000 135.700 ;
    END
  END Y[8]
  PIN Y[9]
    PORT
      LAYER metal1 ;
        RECT 104.400 133.600 106.000 134.400 ;
        RECT 105.300 132.300 105.900 133.600 ;
        RECT 106.800 132.300 107.600 132.400 ;
        RECT 105.300 131.700 107.600 132.300 ;
        RECT 106.800 130.800 107.600 131.700 ;
      LAYER via1 ;
        RECT 105.200 133.600 106.000 134.400 ;
      LAYER metal2 ;
        RECT 105.300 134.400 105.900 144.300 ;
        RECT 105.200 133.600 106.000 134.400 ;
    END
  END Y[9]
  PIN Y[10]
    PORT
      LAYER metal1 ;
        RECT 124.400 28.300 125.200 28.400 ;
        RECT 127.600 28.300 128.400 28.400 ;
        RECT 124.400 28.200 128.400 28.300 ;
        RECT 124.400 27.700 129.200 28.200 ;
        RECT 124.400 27.600 125.200 27.700 ;
        RECT 127.600 27.600 129.200 27.700 ;
        RECT 128.400 27.200 129.200 27.600 ;
        RECT 118.000 24.800 118.800 26.400 ;
        RECT 120.400 13.600 122.000 14.400 ;
      LAYER via1 ;
        RECT 118.000 25.600 118.800 26.400 ;
        RECT 121.200 13.600 122.000 14.400 ;
      LAYER metal2 ;
        RECT 118.000 27.600 118.800 28.400 ;
        RECT 121.200 27.600 122.000 28.400 ;
        RECT 124.400 27.600 125.200 28.400 ;
        RECT 118.100 26.400 118.700 27.600 ;
        RECT 118.000 25.600 118.800 26.400 ;
        RECT 121.300 14.400 121.900 27.600 ;
        RECT 121.200 13.600 122.000 14.400 ;
        RECT 121.300 -2.300 121.900 13.600 ;
      LAYER metal3 ;
        RECT 118.000 28.300 118.800 28.400 ;
        RECT 121.200 28.300 122.000 28.400 ;
        RECT 124.400 28.300 125.200 28.400 ;
        RECT 118.000 27.700 125.200 28.300 ;
        RECT 118.000 27.600 118.800 27.700 ;
        RECT 121.200 27.600 122.000 27.700 ;
        RECT 124.400 27.600 125.200 27.700 ;
    END
  END Y[10]
  PIN Y[11]
    PORT
      LAYER metal1 ;
        RECT 121.200 30.300 122.000 31.200 ;
        RECT 127.600 30.300 128.400 30.400 ;
        RECT 121.200 29.700 128.400 30.300 ;
        RECT 121.200 29.600 122.000 29.700 ;
        RECT 127.600 29.600 128.400 29.700 ;
        RECT 155.600 27.600 157.200 28.400 ;
      LAYER via1 ;
        RECT 156.400 27.600 157.200 28.400 ;
      LAYER metal2 ;
        RECT 127.600 29.600 128.400 30.400 ;
        RECT 127.700 26.400 128.300 29.600 ;
        RECT 156.400 27.600 157.200 28.400 ;
        RECT 156.500 26.400 157.100 27.600 ;
        RECT 127.600 25.600 128.400 26.400 ;
        RECT 156.400 25.600 157.200 26.400 ;
        RECT 156.500 2.400 157.100 25.600 ;
        RECT 151.600 1.600 152.400 2.400 ;
        RECT 156.400 1.600 157.200 2.400 ;
        RECT 151.700 -2.300 152.300 1.600 ;
      LAYER metal3 ;
        RECT 127.600 26.300 128.400 26.400 ;
        RECT 156.400 26.300 157.200 26.400 ;
        RECT 127.600 25.700 157.200 26.300 ;
        RECT 127.600 25.600 128.400 25.700 ;
        RECT 156.400 25.600 157.200 25.700 ;
        RECT 151.600 2.300 152.400 2.400 ;
        RECT 156.400 2.300 157.200 2.400 ;
        RECT 151.600 1.700 157.200 2.300 ;
        RECT 151.600 1.600 152.400 1.700 ;
        RECT 156.400 1.600 157.200 1.700 ;
    END
  END Y[11]
  PIN Y[12]
    PORT
      LAYER metal1 ;
        RECT 95.600 67.600 97.200 68.400 ;
        RECT 106.800 28.200 107.600 28.400 ;
        RECT 106.800 27.600 108.400 28.200 ;
        RECT 107.600 27.200 108.400 27.600 ;
        RECT 95.600 15.600 96.400 17.200 ;
      LAYER metal2 ;
        RECT 95.600 67.600 96.400 68.400 ;
        RECT 95.600 27.600 96.400 28.400 ;
        RECT 106.800 27.600 107.600 28.400 ;
        RECT 95.700 16.400 96.300 27.600 ;
        RECT 95.600 15.600 96.400 16.400 ;
        RECT 95.700 4.400 96.300 15.600 ;
        RECT 95.600 3.600 96.400 4.400 ;
        RECT 100.400 3.600 101.200 4.400 ;
        RECT 100.500 -2.300 101.100 3.600 ;
      LAYER metal3 ;
        RECT 95.600 68.300 96.400 68.400 ;
        RECT 100.400 68.300 101.200 68.400 ;
        RECT 95.600 67.700 101.200 68.300 ;
        RECT 95.600 67.600 96.400 67.700 ;
        RECT 100.400 67.600 101.200 67.700 ;
        RECT 95.600 28.300 96.400 28.400 ;
        RECT 100.400 28.300 101.200 28.400 ;
        RECT 106.800 28.300 107.600 28.400 ;
        RECT 95.600 27.700 107.600 28.300 ;
        RECT 95.600 27.600 96.400 27.700 ;
        RECT 100.400 27.600 101.200 27.700 ;
        RECT 106.800 27.600 107.600 27.700 ;
        RECT 95.600 4.300 96.400 4.400 ;
        RECT 100.400 4.300 101.200 4.400 ;
        RECT 95.600 3.700 101.200 4.300 ;
        RECT 95.600 3.600 96.400 3.700 ;
        RECT 100.400 3.600 101.200 3.700 ;
      LAYER metal4 ;
        RECT 100.200 27.400 101.400 68.600 ;
    END
  END Y[12]
  PIN Y[13]
    PORT
      LAYER metal1 ;
        RECT 100.400 13.600 102.000 14.400 ;
        RECT 98.800 12.300 99.600 12.400 ;
        RECT 100.500 12.300 101.100 13.600 ;
        RECT 103.600 12.300 104.400 12.400 ;
        RECT 98.800 11.700 104.400 12.300 ;
        RECT 98.800 10.800 99.600 11.700 ;
        RECT 103.600 11.600 104.400 11.700 ;
      LAYER metal2 ;
        RECT 103.600 11.600 104.400 12.400 ;
        RECT 103.700 -1.700 104.300 11.600 ;
        RECT 103.700 -2.300 105.900 -1.700 ;
    END
  END Y[13]
  PIN Y[14]
    PORT
      LAYER metal1 ;
        RECT 71.600 24.800 72.400 26.400 ;
        RECT 65.200 15.600 66.000 17.200 ;
      LAYER via1 ;
        RECT 71.600 25.600 72.400 26.400 ;
      LAYER metal2 ;
        RECT 65.200 25.600 66.000 26.400 ;
        RECT 71.600 25.600 72.400 26.400 ;
        RECT 65.300 16.400 65.900 25.600 ;
        RECT 65.200 15.600 66.000 16.400 ;
        RECT 65.300 -2.300 65.900 15.600 ;
      LAYER metal3 ;
        RECT 65.200 26.300 66.000 26.400 ;
        RECT 71.600 26.300 72.400 26.400 ;
        RECT 65.200 25.700 72.400 26.300 ;
        RECT 65.200 25.600 66.000 25.700 ;
        RECT 71.600 25.600 72.400 25.700 ;
    END
  END Y[14]
  PIN Y[15]
    PORT
      LAYER metal1 ;
        RECT 51.600 28.300 53.200 28.400 ;
        RECT 60.400 28.300 61.200 28.400 ;
        RECT 51.600 27.700 61.200 28.300 ;
        RECT 51.600 27.600 53.200 27.700 ;
        RECT 60.400 27.600 61.200 27.700 ;
        RECT 62.000 10.800 62.800 12.400 ;
      LAYER via1 ;
        RECT 62.000 11.600 62.800 12.400 ;
      LAYER metal2 ;
        RECT 60.400 28.300 61.200 28.400 ;
        RECT 60.400 27.700 62.700 28.300 ;
        RECT 60.400 27.600 61.200 27.700 ;
        RECT 62.100 12.400 62.700 27.700 ;
        RECT 62.000 11.600 62.800 12.400 ;
        RECT 62.100 -1.700 62.700 11.600 ;
        RECT 60.500 -2.300 62.700 -1.700 ;
    END
  END Y[15]
  PIN Y[16]
    PORT
      LAYER metal1 ;
        RECT 44.400 55.600 45.200 57.200 ;
        RECT 22.000 53.600 23.600 54.400 ;
        RECT 33.200 50.800 34.000 52.400 ;
      LAYER via1 ;
        RECT 33.200 51.600 34.000 52.400 ;
      LAYER metal2 ;
        RECT 22.000 57.600 22.800 58.400 ;
        RECT 22.100 54.400 22.700 57.600 ;
        RECT 44.400 55.600 45.200 56.400 ;
        RECT 22.000 53.600 22.800 54.400 ;
        RECT 33.200 53.600 34.000 54.400 ;
        RECT 33.300 52.400 33.900 53.600 ;
        RECT 33.200 51.600 34.000 52.400 ;
        RECT 33.300 50.400 33.900 51.600 ;
        RECT 44.500 50.400 45.100 55.600 ;
        RECT 33.200 49.600 34.000 50.400 ;
        RECT 44.400 49.600 45.200 50.400 ;
      LAYER metal3 ;
        RECT 22.000 58.300 22.800 58.400 ;
        RECT -1.900 57.700 22.800 58.300 ;
        RECT 22.000 57.600 22.800 57.700 ;
        RECT 22.000 54.300 22.800 54.400 ;
        RECT 33.200 54.300 34.000 54.400 ;
        RECT 22.000 53.700 34.000 54.300 ;
        RECT 22.000 53.600 22.800 53.700 ;
        RECT 33.200 53.600 34.000 53.700 ;
        RECT 33.200 50.300 34.000 50.400 ;
        RECT 44.400 50.300 45.200 50.400 ;
        RECT 33.200 49.700 45.200 50.300 ;
        RECT 33.200 49.600 34.000 49.700 ;
        RECT 44.400 49.600 45.200 49.700 ;
    END
  END Y[16]
  PIN Y[17]
    PORT
      LAYER metal1 ;
        RECT 36.400 55.600 37.200 57.200 ;
        RECT 59.600 54.400 60.400 54.800 ;
        RECT 58.800 53.800 60.400 54.400 ;
        RECT 58.800 53.600 59.600 53.800 ;
        RECT 32.400 29.600 34.000 30.400 ;
        RECT 36.400 25.600 37.200 26.400 ;
        RECT 36.600 24.800 37.400 25.600 ;
      LAYER via1 ;
        RECT 33.200 29.600 34.000 30.400 ;
      LAYER metal2 ;
        RECT 36.400 55.600 37.200 56.400 ;
        RECT 58.800 55.600 59.600 56.400 ;
        RECT 36.500 30.400 37.100 55.600 ;
        RECT 58.900 54.400 59.500 55.600 ;
        RECT 58.800 53.600 59.600 54.400 ;
        RECT 33.200 29.600 34.000 30.400 ;
        RECT 36.400 29.600 37.200 30.400 ;
        RECT 36.500 26.400 37.100 29.600 ;
        RECT 36.400 25.600 37.200 26.400 ;
        RECT 36.500 -1.700 37.100 25.600 ;
        RECT 36.500 -2.300 38.700 -1.700 ;
      LAYER metal3 ;
        RECT 36.400 56.300 37.200 56.400 ;
        RECT 58.800 56.300 59.600 56.400 ;
        RECT 36.400 55.700 59.600 56.300 ;
        RECT 36.400 55.600 37.200 55.700 ;
        RECT 58.800 55.600 59.600 55.700 ;
        RECT 33.200 30.300 34.000 30.400 ;
        RECT 36.400 30.300 37.200 30.400 ;
        RECT 33.200 29.700 37.200 30.300 ;
        RECT 33.200 29.600 34.000 29.700 ;
        RECT 36.400 29.600 37.200 29.700 ;
    END
  END Y[17]
  PIN Y[18]
    PORT
      LAYER metal1 ;
        RECT 55.600 68.200 56.400 68.400 ;
        RECT 54.800 67.600 56.400 68.200 ;
        RECT 54.800 67.200 55.600 67.600 ;
        RECT 14.000 64.800 14.800 66.400 ;
        RECT 63.600 64.800 64.400 66.400 ;
        RECT 65.200 53.600 66.000 55.200 ;
      LAYER via1 ;
        RECT 55.600 67.600 56.400 68.400 ;
        RECT 14.000 65.600 14.800 66.400 ;
        RECT 63.600 65.600 64.400 66.400 ;
      LAYER metal2 ;
        RECT 55.600 67.600 56.400 68.400 ;
        RECT 55.700 66.400 56.300 67.600 ;
        RECT 14.000 65.600 14.800 66.400 ;
        RECT 55.600 65.600 56.400 66.400 ;
        RECT 63.600 66.300 64.400 66.400 ;
        RECT 63.600 65.700 65.900 66.300 ;
        RECT 63.600 65.600 64.400 65.700 ;
        RECT 65.300 54.400 65.900 65.700 ;
        RECT 65.200 53.600 66.000 54.400 ;
      LAYER metal3 ;
        RECT 14.000 66.300 14.800 66.400 ;
        RECT 55.600 66.300 56.400 66.400 ;
        RECT 63.600 66.300 64.400 66.400 ;
        RECT -1.900 65.700 64.400 66.300 ;
        RECT 14.000 65.600 14.800 65.700 ;
        RECT 55.600 65.600 56.400 65.700 ;
        RECT 63.600 65.600 64.400 65.700 ;
    END
  END Y[18]
  PIN Y[19]
    PORT
      LAYER metal1 ;
        RECT 9.200 70.300 10.000 70.400 ;
        RECT 10.800 70.300 11.600 71.200 ;
        RECT 9.200 69.700 11.600 70.300 ;
        RECT 9.200 69.600 10.000 69.700 ;
        RECT 10.800 69.600 11.600 69.700 ;
        RECT 34.800 67.600 36.400 68.400 ;
      LAYER metal2 ;
        RECT 9.200 69.600 10.000 70.400 ;
        RECT 34.800 69.600 35.600 70.400 ;
        RECT 34.900 68.400 35.500 69.600 ;
        RECT 34.800 67.600 35.600 68.400 ;
      LAYER metal3 ;
        RECT 9.200 70.300 10.000 70.400 ;
        RECT 34.800 70.300 35.600 70.400 ;
        RECT -1.900 69.700 35.600 70.300 ;
        RECT 9.200 69.600 10.000 69.700 ;
        RECT 34.800 69.600 35.600 69.700 ;
    END
  END Y[19]
  PIN Y[20]
    PORT
      LAYER metal1 ;
        RECT 9.200 104.800 10.000 106.400 ;
        RECT 39.600 95.600 40.400 97.200 ;
        RECT 37.200 94.300 38.800 94.400 ;
        RECT 39.700 94.300 40.300 95.600 ;
        RECT 37.200 93.700 40.300 94.300 ;
        RECT 37.200 93.600 38.800 93.700 ;
      LAYER via1 ;
        RECT 9.200 105.600 10.000 106.400 ;
      LAYER metal2 ;
        RECT 9.200 105.600 10.000 106.400 ;
        RECT 9.300 104.400 9.900 105.600 ;
        RECT 9.200 103.600 10.000 104.400 ;
        RECT 9.300 96.400 9.900 103.600 ;
        RECT 9.200 95.600 10.000 96.400 ;
        RECT 39.600 95.600 40.400 96.400 ;
      LAYER metal3 ;
        RECT -1.900 105.700 0.300 106.300 ;
        RECT -0.300 104.300 0.300 105.700 ;
        RECT 9.200 104.300 10.000 104.400 ;
        RECT -0.300 103.700 10.000 104.300 ;
        RECT 9.200 103.600 10.000 103.700 ;
        RECT 9.200 96.300 10.000 96.400 ;
        RECT 39.600 96.300 40.400 96.400 ;
        RECT 9.200 95.700 40.400 96.300 ;
        RECT 9.200 95.600 10.000 95.700 ;
        RECT 39.600 95.600 40.400 95.700 ;
    END
  END Y[20]
  PIN Y[21]
    PORT
      LAYER metal1 ;
        RECT 1.200 95.600 2.000 97.200 ;
        RECT 6.000 92.800 6.800 94.400 ;
      LAYER via1 ;
        RECT 6.000 93.600 6.800 94.400 ;
      LAYER metal2 ;
        RECT 1.200 95.600 2.000 96.400 ;
        RECT 1.300 94.400 1.900 95.600 ;
        RECT 1.200 93.600 2.000 94.400 ;
        RECT 6.000 93.600 6.800 94.400 ;
      LAYER metal3 ;
        RECT 1.200 94.300 2.000 94.400 ;
        RECT 6.000 94.300 6.800 94.400 ;
        RECT -1.900 93.700 6.800 94.300 ;
        RECT 1.200 93.600 2.000 93.700 ;
        RECT 6.000 93.600 6.800 93.700 ;
    END
  END Y[21]
  PIN Y[22]
    PORT
      LAYER metal1 ;
        RECT 8.000 93.800 8.800 94.000 ;
        RECT 7.800 93.200 8.800 93.800 ;
        RECT 7.800 92.400 8.400 93.200 ;
        RECT 4.400 90.800 5.200 92.400 ;
        RECT 7.600 91.600 8.400 92.400 ;
      LAYER via1 ;
        RECT 4.400 91.600 5.200 92.400 ;
      LAYER metal2 ;
        RECT 4.400 91.600 5.200 92.400 ;
        RECT 7.600 91.600 8.400 92.400 ;
        RECT 4.500 90.400 5.100 91.600 ;
        RECT 7.700 90.400 8.300 91.600 ;
        RECT 4.400 89.600 5.200 90.400 ;
        RECT 7.600 89.600 8.400 90.400 ;
      LAYER metal3 ;
        RECT 4.400 90.300 5.200 90.400 ;
        RECT 7.600 90.300 8.400 90.400 ;
        RECT -1.900 89.700 8.400 90.300 ;
        RECT 4.400 89.600 5.200 89.700 ;
        RECT 7.600 89.600 8.400 89.700 ;
    END
  END Y[22]
  PIN Y[23]
    PORT
      LAYER metal1 ;
        RECT 14.800 113.600 15.600 114.400 ;
        RECT 14.800 112.400 15.400 113.600 ;
        RECT 14.000 111.800 15.400 112.400 ;
        RECT 14.000 111.600 14.800 111.800 ;
        RECT 4.400 110.300 5.200 110.400 ;
        RECT 6.000 110.300 6.800 111.200 ;
        RECT 4.400 109.700 6.800 110.300 ;
        RECT 4.400 109.600 5.200 109.700 ;
        RECT 6.000 109.600 6.800 109.700 ;
      LAYER metal2 ;
        RECT 14.000 111.600 14.800 112.400 ;
        RECT 14.100 110.400 14.700 111.600 ;
        RECT 4.400 109.600 5.200 110.400 ;
        RECT 14.000 109.600 14.800 110.400 ;
      LAYER metal3 ;
        RECT 4.400 110.300 5.200 110.400 ;
        RECT 14.000 110.300 14.800 110.400 ;
        RECT -1.900 109.700 14.800 110.300 ;
        RECT 4.400 109.600 5.200 109.700 ;
        RECT 14.000 109.600 14.800 109.700 ;
    END
  END Y[23]
  PIN Y[24]
    PORT
      LAYER metal1 ;
        RECT 22.000 135.600 22.800 137.200 ;
        RECT 16.400 134.400 17.200 134.800 ;
        RECT 16.400 133.800 18.000 134.400 ;
        RECT 17.200 133.600 18.000 133.800 ;
        RECT 26.800 107.600 28.400 108.400 ;
      LAYER metal2 ;
        RECT 22.100 143.700 24.300 144.300 ;
        RECT 22.100 136.400 22.700 143.700 ;
        RECT 22.000 135.600 22.800 136.400 ;
        RECT 22.100 134.400 22.700 135.600 ;
        RECT 17.200 133.600 18.000 134.400 ;
        RECT 22.000 133.600 22.800 134.400 ;
        RECT 26.800 133.600 27.600 134.400 ;
        RECT 26.900 108.400 27.500 133.600 ;
        RECT 26.800 107.600 27.600 108.400 ;
      LAYER metal3 ;
        RECT 17.200 134.300 18.000 134.400 ;
        RECT 22.000 134.300 22.800 134.400 ;
        RECT 26.800 134.300 27.600 134.400 ;
        RECT 17.200 133.700 27.600 134.300 ;
        RECT 17.200 133.600 18.000 133.700 ;
        RECT 22.000 133.600 22.800 133.700 ;
        RECT 26.800 133.600 27.600 133.700 ;
    END
  END Y[24]
  PIN Y[25]
    PORT
      LAYER metal1 ;
        RECT 18.800 130.800 19.600 132.400 ;
        RECT 12.400 130.200 13.200 130.400 ;
        RECT 12.400 129.600 13.800 130.200 ;
        RECT 13.200 128.400 13.800 129.600 ;
        RECT 13.200 127.600 14.000 128.400 ;
      LAYER via1 ;
        RECT 18.800 131.600 19.600 132.400 ;
      LAYER metal2 ;
        RECT 18.900 132.400 19.500 144.300 ;
        RECT 18.800 131.600 19.600 132.400 ;
        RECT 18.900 130.400 19.500 131.600 ;
        RECT 12.400 129.600 13.200 130.400 ;
        RECT 18.800 129.600 19.600 130.400 ;
      LAYER metal3 ;
        RECT 12.400 130.300 13.200 130.400 ;
        RECT 18.800 130.300 19.600 130.400 ;
        RECT 12.400 129.700 19.600 130.300 ;
        RECT 12.400 129.600 13.200 129.700 ;
        RECT 18.800 129.600 19.600 129.700 ;
    END
  END Y[25]
  PIN Y[26]
    PORT
      LAYER metal1 ;
        RECT 39.600 135.600 40.400 137.200 ;
        RECT 63.600 136.300 66.000 136.400 ;
        RECT 68.400 136.300 69.200 137.200 ;
        RECT 63.600 135.700 69.200 136.300 ;
        RECT 63.600 135.600 66.000 135.700 ;
        RECT 68.400 135.600 69.200 135.700 ;
        RECT 34.000 134.400 34.800 134.800 ;
        RECT 33.200 133.800 34.800 134.400 ;
        RECT 33.200 133.600 34.000 133.800 ;
      LAYER via1 ;
        RECT 65.200 135.600 66.000 136.400 ;
      LAYER metal2 ;
        RECT 63.700 136.400 64.300 144.300 ;
        RECT 39.600 135.600 40.400 136.400 ;
        RECT 63.600 135.600 64.400 136.400 ;
        RECT 65.200 135.600 66.000 136.400 ;
        RECT 39.700 134.400 40.300 135.600 ;
        RECT 65.300 134.400 65.900 135.600 ;
        RECT 33.200 133.600 34.000 134.400 ;
        RECT 39.600 133.600 40.400 134.400 ;
        RECT 65.200 133.600 66.000 134.400 ;
      LAYER metal3 ;
        RECT 33.200 134.300 34.000 134.400 ;
        RECT 39.600 134.300 40.400 134.400 ;
        RECT 65.200 134.300 66.000 134.400 ;
        RECT 33.200 133.700 66.000 134.300 ;
        RECT 33.200 133.600 34.000 133.700 ;
        RECT 39.600 133.600 40.400 133.700 ;
        RECT 65.200 133.600 66.000 133.700 ;
    END
  END Y[26]
  PIN Y[27]
    PORT
      LAYER metal1 ;
        RECT 41.200 133.600 42.200 134.400 ;
        RECT 41.600 132.800 42.400 133.600 ;
        RECT 38.000 130.200 38.800 130.400 ;
        RECT 37.400 129.600 38.800 130.200 ;
        RECT 37.400 128.400 38.000 129.600 ;
        RECT 37.200 127.600 38.000 128.400 ;
      LAYER via1 ;
        RECT 38.000 129.600 38.800 130.400 ;
      LAYER metal2 ;
        RECT 41.300 134.400 41.900 144.300 ;
        RECT 41.200 133.600 42.000 134.400 ;
        RECT 41.300 130.400 41.900 133.600 ;
        RECT 38.000 129.600 38.800 130.400 ;
        RECT 41.200 129.600 42.000 130.400 ;
      LAYER metal3 ;
        RECT 38.000 130.300 38.800 130.400 ;
        RECT 41.200 130.300 42.000 130.400 ;
        RECT 38.000 129.700 42.000 130.300 ;
        RECT 38.000 129.600 38.800 129.700 ;
        RECT 41.200 129.600 42.000 129.700 ;
    END
  END Y[27]
  PIN Y[28]
    PORT
      LAYER metal1 ;
        RECT 94.000 135.600 94.800 137.200 ;
        RECT 82.800 109.600 83.600 111.200 ;
        RECT 80.200 96.300 82.000 96.400 ;
        RECT 82.800 96.300 83.600 96.400 ;
        RECT 80.200 95.700 83.600 96.300 ;
        RECT 80.200 95.600 82.000 95.700 ;
        RECT 82.800 95.600 83.600 95.700 ;
      LAYER metal2 ;
        RECT 92.500 136.300 93.100 144.300 ;
        RECT 94.000 136.300 94.800 136.400 ;
        RECT 92.500 135.700 94.800 136.300 ;
        RECT 92.500 120.400 93.100 135.700 ;
        RECT 94.000 135.600 94.800 135.700 ;
        RECT 82.800 119.600 83.600 120.400 ;
        RECT 92.400 119.600 93.200 120.400 ;
        RECT 82.900 110.400 83.500 119.600 ;
        RECT 82.800 109.600 83.600 110.400 ;
        RECT 82.900 96.400 83.500 109.600 ;
        RECT 82.800 95.600 83.600 96.400 ;
      LAYER metal3 ;
        RECT 82.800 120.300 83.600 120.400 ;
        RECT 92.400 120.300 93.200 120.400 ;
        RECT 82.800 119.700 93.200 120.300 ;
        RECT 82.800 119.600 83.600 119.700 ;
        RECT 92.400 119.600 93.200 119.700 ;
    END
  END Y[28]
  PIN Y[29]
    PORT
      LAYER metal1 ;
        RECT 84.400 111.600 85.200 113.200 ;
        RECT 92.400 109.600 93.200 111.200 ;
      LAYER metal2 ;
        RECT 86.100 140.400 86.700 144.300 ;
        RECT 86.000 139.600 86.800 140.400 ;
        RECT 84.400 111.600 85.200 112.400 ;
        RECT 84.500 110.400 85.100 111.600 ;
        RECT 84.400 109.600 85.200 110.400 ;
        RECT 92.400 109.600 93.200 110.400 ;
      LAYER metal3 ;
        RECT 84.400 140.300 85.200 140.400 ;
        RECT 86.000 140.300 86.800 140.400 ;
        RECT 84.400 139.700 86.800 140.300 ;
        RECT 84.400 139.600 85.200 139.700 ;
        RECT 86.000 139.600 86.800 139.700 ;
        RECT 84.400 110.300 85.200 110.400 ;
        RECT 92.400 110.300 93.200 110.400 ;
        RECT 84.400 109.700 93.200 110.300 ;
        RECT 84.400 109.600 85.200 109.700 ;
        RECT 92.400 109.600 93.200 109.700 ;
      LAYER metal4 ;
        RECT 84.200 109.400 85.400 140.600 ;
    END
  END Y[29]
  PIN Y[30]
    PORT
      LAYER metal1 ;
        RECT 87.600 108.300 88.400 108.400 ;
        RECT 89.200 108.300 90.000 108.400 ;
        RECT 87.600 107.700 90.000 108.300 ;
        RECT 87.600 106.800 88.400 107.700 ;
        RECT 89.200 107.600 90.000 107.700 ;
        RECT 89.300 106.400 89.900 107.600 ;
        RECT 89.200 104.800 90.000 106.400 ;
      LAYER metal2 ;
        RECT 89.300 108.400 89.900 144.300 ;
        RECT 89.200 107.600 90.000 108.400 ;
    END
  END Y[30]
  PIN Y[31]
    PORT
      LAYER metal1 ;
        RECT 116.400 70.300 117.200 70.400 ;
        RECT 118.000 70.300 118.800 70.400 ;
        RECT 116.400 69.700 118.800 70.300 ;
        RECT 116.400 68.800 117.200 69.700 ;
        RECT 118.000 68.800 118.800 69.700 ;
        RECT 122.800 68.800 123.600 70.400 ;
        RECT 135.600 68.800 136.400 70.400 ;
      LAYER via1 ;
        RECT 118.000 69.600 118.800 70.400 ;
        RECT 122.800 69.600 123.600 70.400 ;
        RECT 135.600 69.600 136.400 70.400 ;
      LAYER metal2 ;
        RECT 118.000 69.600 118.800 70.400 ;
        RECT 122.800 69.600 123.600 70.400 ;
        RECT 135.600 69.600 136.400 70.400 ;
      LAYER metal3 ;
        RECT 118.000 70.300 118.800 70.400 ;
        RECT 122.800 70.300 123.600 70.400 ;
        RECT 135.600 70.300 136.400 70.400 ;
        RECT 118.000 69.700 182.700 70.300 ;
        RECT 118.000 69.600 118.800 69.700 ;
        RECT 122.800 69.600 123.600 69.700 ;
        RECT 135.600 69.600 136.400 69.700 ;
    END
  END Y[31]
  PIN O[0]
    PORT
      LAYER metal1 ;
        RECT 150.000 132.400 150.800 139.800 ;
        RECT 150.200 130.200 150.800 132.400 ;
        RECT 150.000 122.200 150.800 130.200 ;
      LAYER via1 ;
        RECT 150.000 137.600 150.800 138.400 ;
      LAYER metal2 ;
        RECT 148.500 143.700 150.700 144.300 ;
        RECT 150.100 138.400 150.700 143.700 ;
        RECT 150.000 137.600 150.800 138.400 ;
    END
  END O[0]
  PIN O[1]
    PORT
      LAYER metal1 ;
        RECT 169.200 111.800 170.000 119.800 ;
        RECT 169.400 109.600 170.000 111.800 ;
        RECT 169.200 102.200 170.000 109.600 ;
      LAYER via1 ;
        RECT 169.200 115.600 170.000 116.400 ;
      LAYER metal2 ;
        RECT 169.200 115.600 170.000 116.400 ;
      LAYER metal3 ;
        RECT 169.200 116.300 170.000 116.400 ;
        RECT 169.200 115.700 182.700 116.300 ;
        RECT 169.200 115.600 170.000 115.700 ;
    END
  END O[1]
  PIN O[2]
    PORT
      LAYER metal1 ;
        RECT 148.400 12.400 149.200 19.800 ;
        RECT 148.600 10.200 149.200 12.400 ;
        RECT 148.400 2.200 149.200 10.200 ;
      LAYER via1 ;
        RECT 148.400 3.600 149.200 4.400 ;
      LAYER metal2 ;
        RECT 148.400 3.600 149.200 4.400 ;
        RECT 148.500 -1.700 149.100 3.600 ;
        RECT 146.900 -2.300 149.100 -1.700 ;
    END
  END O[2]
  PIN O[3]
    PORT
      LAYER metal1 ;
        RECT 172.400 54.300 173.200 59.800 ;
        RECT 174.000 54.300 174.800 54.400 ;
        RECT 172.400 53.700 174.800 54.300 ;
        RECT 172.400 52.400 173.200 53.700 ;
        RECT 174.000 53.600 174.800 53.700 ;
        RECT 172.600 50.200 173.200 52.400 ;
        RECT 172.400 42.200 173.200 50.200 ;
      LAYER metal2 ;
        RECT 174.000 53.600 174.800 54.400 ;
      LAYER metal3 ;
        RECT 174.000 54.300 174.800 54.400 ;
        RECT 174.000 53.700 182.700 54.300 ;
        RECT 174.000 53.600 174.800 53.700 ;
    END
  END O[3]
  PIN O[4]
    PORT
      LAYER metal1 ;
        RECT 140.400 132.400 141.200 139.800 ;
        RECT 140.600 130.200 141.200 132.400 ;
        RECT 140.400 122.200 141.200 130.200 ;
      LAYER via1 ;
        RECT 140.400 137.600 141.200 138.400 ;
      LAYER metal2 ;
        RECT 137.300 140.400 137.900 144.300 ;
        RECT 137.200 139.600 138.000 140.400 ;
        RECT 140.400 139.600 141.200 140.400 ;
        RECT 140.500 138.400 141.100 139.600 ;
        RECT 140.400 137.600 141.200 138.400 ;
      LAYER metal3 ;
        RECT 137.200 140.300 138.000 140.400 ;
        RECT 140.400 140.300 141.200 140.400 ;
        RECT 137.200 139.700 141.200 140.300 ;
        RECT 137.200 139.600 138.000 139.700 ;
        RECT 140.400 139.600 141.200 139.700 ;
    END
  END O[4]
  PIN O[5]
    PORT
      LAYER metal1 ;
        RECT 135.600 132.400 136.400 139.800 ;
        RECT 135.800 130.200 136.400 132.400 ;
        RECT 135.600 122.200 136.400 130.200 ;
      LAYER via1 ;
        RECT 135.600 137.600 136.400 138.400 ;
      LAYER metal2 ;
        RECT 132.500 140.400 133.100 144.300 ;
        RECT 132.400 139.600 133.200 140.400 ;
        RECT 135.600 139.600 136.400 140.400 ;
        RECT 135.700 138.400 136.300 139.600 ;
        RECT 135.600 137.600 136.400 138.400 ;
      LAYER metal3 ;
        RECT 132.400 140.300 133.200 140.400 ;
        RECT 135.600 140.300 136.400 140.400 ;
        RECT 132.400 139.700 136.400 140.300 ;
        RECT 132.400 139.600 133.200 139.700 ;
        RECT 135.600 139.600 136.400 139.700 ;
    END
  END O[5]
  PIN O[6]
    PORT
      LAYER metal1 ;
        RECT 143.600 12.400 144.400 19.800 ;
        RECT 143.800 10.200 144.400 12.400 ;
        RECT 143.600 2.200 144.400 10.200 ;
      LAYER via1 ;
        RECT 143.600 3.600 144.400 4.400 ;
      LAYER metal2 ;
        RECT 143.600 3.600 144.400 4.400 ;
        RECT 143.700 2.400 144.300 3.600 ;
        RECT 140.400 1.600 141.200 2.400 ;
        RECT 143.600 1.600 144.400 2.400 ;
        RECT 140.500 -2.300 141.100 1.600 ;
      LAYER metal3 ;
        RECT 140.400 2.300 141.200 2.400 ;
        RECT 143.600 2.300 144.400 2.400 ;
        RECT 140.400 1.700 144.400 2.300 ;
        RECT 140.400 1.600 141.200 1.700 ;
        RECT 143.600 1.600 144.400 1.700 ;
    END
  END O[6]
  PIN O[7]
    PORT
      LAYER metal1 ;
        RECT 174.000 12.400 174.800 19.800 ;
        RECT 174.000 10.200 174.600 12.400 ;
        RECT 174.000 2.200 174.800 10.200 ;
      LAYER via1 ;
        RECT 174.000 3.600 174.800 4.400 ;
      LAYER metal2 ;
        RECT 174.000 3.600 174.800 4.400 ;
        RECT 174.100 -1.700 174.700 3.600 ;
        RECT 174.100 -2.300 176.300 -1.700 ;
    END
  END O[7]
  PIN O[8]
    PORT
      LAYER metal1 ;
        RECT 92.400 31.800 93.200 39.800 ;
        RECT 92.400 29.600 93.000 31.800 ;
        RECT 92.400 22.200 93.200 29.600 ;
      LAYER via1 ;
        RECT 92.400 23.600 93.200 24.400 ;
      LAYER metal2 ;
        RECT 92.400 23.600 93.200 24.400 ;
        RECT 92.500 -1.700 93.100 23.600 ;
        RECT 92.500 -2.300 94.700 -1.700 ;
    END
  END O[8]
  PIN O[9]
    PORT
      LAYER metal1 ;
        RECT 166.000 12.400 166.800 19.800 ;
        RECT 166.200 10.200 166.800 12.400 ;
        RECT 166.000 2.200 166.800 10.200 ;
      LAYER via1 ;
        RECT 166.000 3.600 166.800 4.400 ;
      LAYER metal2 ;
        RECT 166.000 3.600 166.800 4.400 ;
        RECT 166.100 -1.700 166.700 3.600 ;
        RECT 164.500 -2.300 166.700 -1.700 ;
    END
  END O[9]
  PIN O[10]
    PORT
      LAYER metal1 ;
        RECT 94.000 12.400 94.800 19.800 ;
        RECT 94.200 10.200 94.800 12.400 ;
        RECT 94.000 2.200 94.800 10.200 ;
      LAYER via1 ;
        RECT 94.000 3.600 94.800 4.400 ;
      LAYER metal2 ;
        RECT 94.000 3.600 94.800 4.400 ;
        RECT 94.100 2.400 94.700 3.600 ;
        RECT 94.000 1.600 94.800 2.400 ;
        RECT 97.200 1.600 98.000 2.400 ;
        RECT 97.300 -2.300 97.900 1.600 ;
      LAYER metal3 ;
        RECT 94.000 2.300 94.800 2.400 ;
        RECT 97.200 2.300 98.000 2.400 ;
        RECT 94.000 1.700 98.000 2.300 ;
        RECT 94.000 1.600 94.800 1.700 ;
        RECT 97.200 1.600 98.000 1.700 ;
    END
  END O[10]
  PIN O[11]
    PORT
      LAYER metal1 ;
        RECT 34.800 12.400 35.600 19.800 ;
        RECT 34.800 10.200 35.400 12.400 ;
        RECT 34.800 2.200 35.600 10.200 ;
      LAYER via1 ;
        RECT 34.800 3.600 35.600 4.400 ;
      LAYER metal2 ;
        RECT 34.800 3.600 35.600 4.400 ;
        RECT 34.900 -2.300 35.500 3.600 ;
    END
  END O[11]
  PIN O[12]
    PORT
      LAYER metal1 ;
        RECT 1.200 12.400 2.000 19.800 ;
        RECT 1.200 10.200 1.800 12.400 ;
        RECT 1.200 2.200 2.000 10.200 ;
      LAYER via1 ;
        RECT 1.200 7.600 2.000 8.400 ;
      LAYER metal2 ;
        RECT 1.200 9.600 2.000 10.400 ;
        RECT 1.300 8.400 1.900 9.600 ;
        RECT 1.200 7.600 2.000 8.400 ;
      LAYER metal3 ;
        RECT 1.200 10.300 2.000 10.400 ;
        RECT -1.900 9.700 2.000 10.300 ;
        RECT 1.200 9.600 2.000 9.700 ;
    END
  END O[12]
  PIN O[13]
    PORT
      LAYER metal1 ;
        RECT 17.200 12.400 18.000 19.800 ;
        RECT 17.200 10.200 17.800 12.400 ;
        RECT 17.200 2.200 18.000 10.200 ;
      LAYER via1 ;
        RECT 17.200 3.600 18.000 4.400 ;
      LAYER metal2 ;
        RECT 17.200 3.600 18.000 4.400 ;
        RECT 17.300 -1.700 17.900 3.600 ;
        RECT 17.300 -2.300 19.500 -1.700 ;
    END
  END O[13]
  PIN O[14]
    PORT
      LAYER metal1 ;
        RECT 60.400 12.400 61.200 19.800 ;
        RECT 60.600 10.200 61.200 12.400 ;
        RECT 60.400 2.200 61.200 10.200 ;
      LAYER via1 ;
        RECT 60.400 3.600 61.200 4.400 ;
      LAYER metal2 ;
        RECT 60.400 3.600 61.200 4.400 ;
        RECT 60.500 2.400 61.100 3.600 ;
        RECT 57.200 1.600 58.000 2.400 ;
        RECT 60.400 1.600 61.200 2.400 ;
        RECT 57.300 -2.300 57.900 1.600 ;
      LAYER metal3 ;
        RECT 57.200 2.300 58.000 2.400 ;
        RECT 60.400 2.300 61.200 2.400 ;
        RECT 57.200 1.700 61.200 2.300 ;
        RECT 57.200 1.600 58.000 1.700 ;
        RECT 60.400 1.600 61.200 1.700 ;
    END
  END O[14]
  PIN O[15]
    PORT
      LAYER metal1 ;
        RECT 167.600 52.400 168.400 59.800 ;
        RECT 167.800 50.200 168.400 52.400 ;
        RECT 167.600 42.200 168.400 50.200 ;
      LAYER via1 ;
        RECT 167.600 47.600 168.400 48.400 ;
      LAYER metal2 ;
        RECT 167.600 47.600 168.400 48.400 ;
      LAYER metal3 ;
        RECT 167.600 48.300 168.400 48.400 ;
        RECT 182.100 48.300 182.700 50.300 ;
        RECT 167.600 47.700 182.700 48.300 ;
        RECT 167.600 47.600 168.400 47.700 ;
    END
  END O[15]
  PIN O[16]
    PORT
      LAYER metal1 ;
        RECT 6.000 12.400 6.800 19.800 ;
        RECT 6.000 10.200 6.600 12.400 ;
        RECT 6.000 2.200 6.800 10.200 ;
      LAYER via1 ;
        RECT 6.000 13.600 6.800 14.400 ;
      LAYER metal2 ;
        RECT 6.000 13.600 6.800 14.400 ;
      LAYER metal3 ;
        RECT 6.000 14.300 6.800 14.400 ;
        RECT -1.900 13.700 6.800 14.300 ;
        RECT 6.000 13.600 6.800 13.700 ;
    END
  END O[16]
  PIN O[17]
    PORT
      LAYER metal1 ;
        RECT 177.200 98.300 178.000 99.800 ;
        RECT 178.800 98.300 179.600 98.400 ;
        RECT 177.200 97.700 179.600 98.300 ;
        RECT 177.200 92.400 178.000 97.700 ;
        RECT 178.800 97.600 179.600 97.700 ;
        RECT 177.400 90.200 178.000 92.400 ;
        RECT 177.200 82.200 178.000 90.200 ;
      LAYER metal2 ;
        RECT 178.800 101.600 179.600 102.400 ;
        RECT 178.900 98.400 179.500 101.600 ;
        RECT 178.800 97.600 179.600 98.400 ;
      LAYER metal3 ;
        RECT 178.800 102.300 179.600 102.400 ;
        RECT 178.800 101.700 182.700 102.300 ;
        RECT 178.800 101.600 179.600 101.700 ;
    END
  END O[17]
  PIN O[18]
    PORT
      LAYER metal1 ;
        RECT 159.600 132.400 160.400 139.800 ;
        RECT 159.800 130.200 160.400 132.400 ;
        RECT 159.600 122.200 160.400 130.200 ;
      LAYER via1 ;
        RECT 159.600 137.600 160.400 138.400 ;
      LAYER metal2 ;
        RECT 158.100 143.700 160.300 144.300 ;
        RECT 159.700 138.400 160.300 143.700 ;
        RECT 159.600 137.600 160.400 138.400 ;
    END
  END O[18]
  PIN O[19]
    PORT
      LAYER metal1 ;
        RECT 1.200 132.400 2.000 139.800 ;
        RECT 1.200 130.200 1.800 132.400 ;
        RECT 1.200 122.200 2.000 130.200 ;
      LAYER via1 ;
        RECT 1.200 127.600 2.000 128.400 ;
      LAYER metal2 ;
        RECT 1.200 129.600 2.000 130.400 ;
        RECT 1.300 128.400 1.900 129.600 ;
        RECT 1.200 127.600 2.000 128.400 ;
      LAYER metal3 ;
        RECT 1.200 130.300 2.000 130.400 ;
        RECT -1.900 129.700 2.000 130.300 ;
        RECT 1.200 129.600 2.000 129.700 ;
    END
  END O[19]
  PIN O[20]
    PORT
      LAYER metal1 ;
        RECT 174.000 31.800 174.800 39.800 ;
        RECT 174.200 29.600 174.800 31.800 ;
        RECT 174.000 28.300 174.800 29.600 ;
        RECT 178.800 28.300 179.600 28.400 ;
        RECT 174.000 27.700 179.600 28.300 ;
        RECT 174.000 22.200 174.800 27.700 ;
        RECT 178.800 27.600 179.600 27.700 ;
      LAYER metal2 ;
        RECT 178.800 29.600 179.600 30.400 ;
        RECT 178.900 28.400 179.500 29.600 ;
        RECT 178.800 27.600 179.600 28.400 ;
      LAYER metal3 ;
        RECT 178.800 30.300 179.600 30.400 ;
        RECT 178.800 29.700 182.700 30.300 ;
        RECT 178.800 29.600 179.600 29.700 ;
    END
  END O[20]
  PIN O[21]
    PORT
      LAYER metal1 ;
        RECT 164.400 71.800 165.200 79.800 ;
        RECT 164.400 69.600 165.000 71.800 ;
        RECT 164.400 62.200 165.200 69.600 ;
      LAYER via1 ;
        RECT 164.400 77.600 165.200 78.400 ;
      LAYER metal2 ;
        RECT 164.400 87.600 165.200 88.400 ;
        RECT 164.500 78.400 165.100 87.600 ;
        RECT 164.400 77.600 165.200 78.400 ;
      LAYER metal3 ;
        RECT 164.400 88.300 165.200 88.400 ;
        RECT 182.100 88.300 182.700 90.300 ;
        RECT 164.400 87.700 182.700 88.300 ;
        RECT 164.400 87.600 165.200 87.700 ;
    END
  END O[21]
  PIN O[22]
    PORT
      LAYER metal1 ;
        RECT 1.200 52.400 2.000 59.800 ;
        RECT 1.200 50.200 1.800 52.400 ;
        RECT 1.200 42.200 2.000 50.200 ;
      LAYER via1 ;
        RECT 1.200 47.600 2.000 48.400 ;
      LAYER metal2 ;
        RECT 1.200 49.600 2.000 50.400 ;
        RECT 1.300 48.400 1.900 49.600 ;
        RECT 1.200 47.600 2.000 48.400 ;
      LAYER metal3 ;
        RECT 1.200 50.300 2.000 50.400 ;
        RECT -1.900 49.700 2.000 50.300 ;
        RECT 1.200 49.600 2.000 49.700 ;
    END
  END O[22]
  PIN O[23]
    PORT
      LAYER metal1 ;
        RECT 6.000 52.400 6.800 59.800 ;
        RECT 6.000 50.200 6.600 52.400 ;
        RECT 6.000 42.200 6.800 50.200 ;
      LAYER via1 ;
        RECT 6.000 53.600 6.800 54.400 ;
      LAYER metal2 ;
        RECT 6.000 53.600 6.800 54.400 ;
      LAYER metal3 ;
        RECT 6.000 54.300 6.800 54.400 ;
        RECT -1.900 53.700 6.800 54.300 ;
        RECT 6.000 53.600 6.800 53.700 ;
    END
  END O[23]
  PIN O[24]
    PORT
      LAYER metal1 ;
        RECT 177.200 71.800 178.000 79.800 ;
        RECT 177.400 69.600 178.000 71.800 ;
        RECT 177.200 62.200 178.000 69.600 ;
      LAYER via1 ;
        RECT 177.200 77.600 178.000 78.400 ;
      LAYER metal2 ;
        RECT 177.200 81.600 178.000 82.400 ;
        RECT 177.300 78.400 177.900 81.600 ;
        RECT 177.200 77.600 178.000 78.400 ;
      LAYER metal3 ;
        RECT 177.200 82.300 178.000 82.400 ;
        RECT 177.200 81.700 182.700 82.300 ;
        RECT 177.200 81.600 178.000 81.700 ;
    END
  END O[24]
  PIN O[25]
    PORT
      LAYER metal1 ;
        RECT 154.800 132.400 155.600 139.800 ;
        RECT 155.000 130.200 155.600 132.400 ;
        RECT 154.800 122.200 155.600 130.200 ;
      LAYER via1 ;
        RECT 154.800 137.600 155.600 138.400 ;
      LAYER metal2 ;
        RECT 153.300 143.700 155.500 144.300 ;
        RECT 154.900 138.400 155.500 143.700 ;
        RECT 154.800 137.600 155.600 138.400 ;
    END
  END O[25]
  PIN O[26]
    PORT
      LAYER metal1 ;
        RECT 172.400 71.800 173.200 79.800 ;
        RECT 172.600 69.600 173.200 71.800 ;
        RECT 172.400 62.200 173.200 69.600 ;
      LAYER via1 ;
        RECT 172.400 77.600 173.200 78.400 ;
      LAYER metal2 ;
        RECT 172.400 79.600 173.200 80.400 ;
        RECT 172.500 78.400 173.100 79.600 ;
        RECT 172.400 77.600 173.200 78.400 ;
      LAYER metal3 ;
        RECT 177.200 84.300 178.000 84.400 ;
        RECT 182.100 84.300 182.700 86.300 ;
        RECT 177.200 83.700 182.700 84.300 ;
        RECT 177.200 83.600 178.000 83.700 ;
        RECT 172.400 80.300 173.200 80.400 ;
        RECT 177.200 80.300 178.000 80.400 ;
        RECT 172.400 79.700 178.000 80.300 ;
        RECT 172.400 79.600 173.200 79.700 ;
        RECT 177.200 79.600 178.000 79.700 ;
      LAYER metal4 ;
        RECT 177.000 79.400 178.200 84.600 ;
    END
  END O[26]
  PIN O[27]
    PORT
      LAYER metal1 ;
        RECT 1.200 71.800 2.000 79.800 ;
        RECT 1.200 69.600 1.800 71.800 ;
        RECT 1.200 62.200 2.000 69.600 ;
      LAYER via1 ;
        RECT 1.200 73.600 2.000 74.400 ;
      LAYER metal2 ;
        RECT 1.200 73.600 2.000 74.400 ;
      LAYER metal3 ;
        RECT 1.200 74.300 2.000 74.400 ;
        RECT -1.900 73.700 2.000 74.300 ;
        RECT 1.200 73.600 2.000 73.700 ;
    END
  END O[27]
  PIN O[28]
    PORT
      LAYER metal1 ;
        RECT 164.400 132.400 165.200 139.800 ;
        RECT 164.600 130.200 165.200 132.400 ;
        RECT 164.400 122.200 165.200 130.200 ;
      LAYER via1 ;
        RECT 164.400 137.600 165.200 138.400 ;
      LAYER metal2 ;
        RECT 162.900 143.700 165.100 144.300 ;
        RECT 164.500 138.400 165.100 143.700 ;
        RECT 164.400 137.600 165.200 138.400 ;
    END
  END O[28]
  PIN O[29]
    PORT
      LAYER metal1 ;
        RECT 174.000 132.400 174.800 139.800 ;
        RECT 174.200 130.200 174.800 132.400 ;
        RECT 174.000 122.200 174.800 130.200 ;
      LAYER via1 ;
        RECT 174.000 137.600 174.800 138.400 ;
      LAYER metal2 ;
        RECT 172.500 143.700 174.700 144.300 ;
        RECT 174.100 138.400 174.700 143.700 ;
        RECT 174.000 137.600 174.800 138.400 ;
    END
  END O[29]
  PIN O[30]
    PORT
      LAYER metal1 ;
        RECT 145.200 132.400 146.000 139.800 ;
        RECT 145.400 130.200 146.000 132.400 ;
        RECT 145.200 122.200 146.000 130.200 ;
      LAYER via1 ;
        RECT 145.200 137.600 146.000 138.400 ;
      LAYER metal2 ;
        RECT 142.100 140.400 142.700 144.300 ;
        RECT 142.000 139.600 142.800 140.400 ;
        RECT 145.200 139.600 146.000 140.400 ;
        RECT 145.300 138.400 145.900 139.600 ;
        RECT 145.200 137.600 146.000 138.400 ;
      LAYER metal3 ;
        RECT 142.000 140.300 142.800 140.400 ;
        RECT 145.200 140.300 146.000 140.400 ;
        RECT 142.000 139.700 146.000 140.300 ;
        RECT 142.000 139.600 142.800 139.700 ;
        RECT 145.200 139.600 146.000 139.700 ;
    END
  END O[30]
  PIN O[31]
    PORT
      LAYER metal1 ;
        RECT 169.200 132.400 170.000 139.800 ;
        RECT 169.400 130.200 170.000 132.400 ;
        RECT 169.200 122.200 170.000 130.200 ;
      LAYER via1 ;
        RECT 169.200 137.600 170.000 138.400 ;
      LAYER metal2 ;
        RECT 167.700 143.700 169.900 144.300 ;
        RECT 169.300 138.400 169.900 143.700 ;
        RECT 169.200 137.600 170.000 138.400 ;
    END
  END O[31]
  OBS
      LAYER metal1 ;
        RECT 4.400 135.200 5.200 139.800 ;
        RECT 6.600 136.800 7.400 139.800 ;
        RECT 3.000 134.600 5.200 135.200 ;
        RECT 6.000 135.800 7.400 136.800 ;
        RECT 10.800 135.800 11.600 139.800 ;
        RECT 12.400 135.800 13.200 139.800 ;
        RECT 14.000 136.000 14.800 139.800 ;
        RECT 17.200 136.000 18.000 139.800 ;
        RECT 14.000 135.800 18.000 136.000 ;
        RECT 20.400 137.800 21.200 139.800 ;
        RECT 20.400 136.400 21.000 137.800 ;
        RECT 3.000 131.600 3.600 134.600 ;
        RECT 2.400 130.800 3.600 131.600 ;
        RECT 3.000 130.200 3.600 130.800 ;
        RECT 6.000 132.400 6.600 135.800 ;
        RECT 10.800 135.600 11.400 135.800 ;
        RECT 9.600 135.200 11.400 135.600 ;
        RECT 7.200 135.000 11.400 135.200 ;
        RECT 7.200 134.600 10.200 135.000 ;
        RECT 7.200 134.400 8.000 134.600 ;
        RECT 12.600 134.400 13.200 135.800 ;
        RECT 14.200 135.400 17.800 135.800 ;
        RECT 20.400 135.600 21.200 136.400 ;
        RECT 23.600 135.800 24.400 139.800 ;
        RECT 26.800 137.800 27.600 139.800 ;
        RECT 20.400 134.400 21.000 135.600 ;
        RECT 6.000 131.600 6.800 132.400 ;
        RECT 6.000 130.200 6.600 131.600 ;
        RECT 7.400 131.000 8.000 134.400 ;
        RECT 8.800 133.800 9.600 134.000 ;
        RECT 8.800 133.200 9.800 133.800 ;
        RECT 9.200 132.400 9.800 133.200 ;
        RECT 10.800 132.800 11.600 134.400 ;
        RECT 12.400 133.600 15.000 134.400 ;
        RECT 9.200 131.600 10.000 132.400 ;
        RECT 12.400 132.300 13.200 132.400 ;
        RECT 14.400 132.300 15.000 133.600 ;
        RECT 20.400 133.600 21.200 134.400 ;
        RECT 12.400 131.700 15.000 132.300 ;
        RECT 12.400 131.600 13.200 131.700 ;
        RECT 7.400 130.400 9.800 131.000 ;
        RECT 3.000 129.600 5.200 130.200 ;
        RECT 4.400 122.200 5.200 129.600 ;
        RECT 6.000 122.200 6.800 130.200 ;
        RECT 9.200 126.200 9.800 130.400 ;
        RECT 14.400 130.200 15.000 131.700 ;
        RECT 15.600 132.300 16.400 133.200 ;
        RECT 17.200 132.300 18.000 132.400 ;
        RECT 15.600 131.700 18.000 132.300 ;
        RECT 15.600 131.600 16.400 131.700 ;
        RECT 17.200 131.600 18.000 131.700 ;
        RECT 20.400 130.200 21.000 133.600 ;
        RECT 23.600 132.400 24.200 135.800 ;
        RECT 26.800 135.600 27.400 137.800 ;
        RECT 28.400 135.600 29.200 137.200 ;
        RECT 30.000 135.600 30.800 137.200 ;
        RECT 25.000 135.000 27.400 135.600 ;
        RECT 23.600 131.600 24.400 132.400 ;
        RECT 25.000 132.000 25.600 135.000 ;
        RECT 26.600 134.300 27.600 134.400 ;
        RECT 31.600 134.300 32.400 139.800 ;
        RECT 33.200 136.000 34.000 139.800 ;
        RECT 36.400 136.000 37.200 139.800 ;
        RECT 33.200 135.800 37.200 136.000 ;
        RECT 38.000 135.800 38.800 139.800 ;
        RECT 41.200 137.800 42.000 139.800 ;
        RECT 33.400 135.400 37.000 135.800 ;
        RECT 38.000 134.400 38.600 135.800 ;
        RECT 41.400 135.600 42.000 137.800 ;
        RECT 44.400 136.300 45.200 139.800 ;
        RECT 47.600 137.800 48.400 139.800 ;
        RECT 60.400 137.800 61.200 139.800 ;
        RECT 63.600 138.400 64.400 139.800 ;
        RECT 46.000 136.300 46.800 137.200 ;
        RECT 44.400 135.800 46.800 136.300 ;
        RECT 44.500 135.700 46.800 135.800 ;
        RECT 41.400 135.000 43.800 135.600 ;
        RECT 26.600 133.700 32.400 134.300 ;
        RECT 26.600 133.600 27.600 133.700 ;
        RECT 26.400 132.800 27.200 133.600 ;
        RECT 31.600 132.300 32.400 133.700 ;
        RECT 36.200 133.600 38.800 134.400 ;
        RECT 33.200 132.300 34.000 132.400 ;
        RECT 23.600 130.400 24.200 131.600 ;
        RECT 25.000 131.400 25.800 132.000 ;
        RECT 31.600 131.700 34.000 132.300 ;
        RECT 25.000 131.200 29.200 131.400 ;
        RECT 25.200 130.800 29.200 131.200 ;
        RECT 23.600 130.200 24.400 130.400 ;
        RECT 14.400 129.600 15.400 130.200 ;
        RECT 9.200 122.200 10.000 126.200 ;
        RECT 14.600 122.200 15.400 129.600 ;
        RECT 19.400 129.400 21.200 130.200 ;
        RECT 23.600 129.600 25.000 130.200 ;
        RECT 19.400 122.200 20.200 129.400 ;
        RECT 24.200 122.200 25.000 129.600 ;
        RECT 28.400 122.200 29.200 130.800 ;
        RECT 31.600 122.200 32.400 131.700 ;
        RECT 33.200 131.600 34.000 131.700 ;
        RECT 34.800 131.600 35.600 133.200 ;
        RECT 36.200 130.200 36.800 133.600 ;
        RECT 43.200 132.000 43.800 135.000 ;
        RECT 44.600 132.400 45.200 135.700 ;
        RECT 46.000 135.600 46.800 135.700 ;
        RECT 47.800 134.400 48.400 137.800 ;
        RECT 60.000 137.600 61.200 137.800 ;
        RECT 63.400 137.800 64.400 138.400 ;
        RECT 63.400 137.600 64.000 137.800 ;
        RECT 60.000 137.000 64.000 137.600 ;
        RECT 60.000 134.400 60.600 137.000 ;
        RECT 70.000 136.300 70.800 139.800 ;
        RECT 71.800 136.400 72.600 137.200 ;
        RECT 71.600 136.300 72.400 136.400 ;
        RECT 70.000 135.700 72.400 136.300 ;
        RECT 73.200 135.800 74.000 139.800 ;
        RECT 78.000 136.000 78.800 139.800 ;
        RECT 81.200 139.200 85.200 139.800 ;
        RECT 81.200 136.000 82.000 139.200 ;
        RECT 78.000 135.800 82.000 136.000 ;
        RECT 82.800 135.800 83.600 138.600 ;
        RECT 84.400 135.800 85.200 139.200 ;
        RECT 89.200 135.800 90.000 139.800 ;
        RECT 90.600 136.400 91.400 137.200 ;
        RECT 90.800 136.300 91.600 136.400 ;
        RECT 92.400 136.300 93.200 139.800 ;
        RECT 47.600 134.300 48.400 134.400 ;
        RECT 57.200 134.300 58.000 134.400 ;
        RECT 47.600 133.700 58.000 134.300 ;
        RECT 47.600 133.600 48.400 133.700 ;
        RECT 57.200 133.600 58.000 133.700 ;
        RECT 60.000 133.600 61.200 134.400 ;
        RECT 62.800 133.600 64.400 134.400 ;
        RECT 43.000 131.400 43.800 132.000 ;
        RECT 44.400 131.600 45.200 132.400 ;
        RECT 35.800 129.600 36.800 130.200 ;
        RECT 39.600 131.200 43.800 131.400 ;
        RECT 39.600 130.800 43.600 131.200 ;
        RECT 35.800 124.400 36.600 129.600 ;
        RECT 34.800 123.600 36.600 124.400 ;
        RECT 35.800 122.200 36.600 123.600 ;
        RECT 39.600 122.200 40.400 130.800 ;
        RECT 44.600 130.200 45.200 131.600 ;
        RECT 47.800 130.200 48.400 133.600 ;
        RECT 49.200 130.800 50.000 132.400 ;
        RECT 60.000 130.400 60.600 133.600 ;
        RECT 61.200 131.600 62.800 132.400 ;
        RECT 43.800 129.600 45.200 130.200 ;
        RECT 43.800 122.200 44.600 129.600 ;
        RECT 47.600 129.400 49.400 130.200 ;
        RECT 57.200 129.800 60.600 130.400 ;
        RECT 57.200 129.600 58.000 129.800 ;
        RECT 48.600 122.200 49.400 129.400 ;
        RECT 57.400 129.000 58.000 129.600 ;
        RECT 59.000 129.000 62.600 129.200 ;
        RECT 55.600 123.000 56.400 129.000 ;
        RECT 57.200 123.400 58.000 129.000 ;
        RECT 58.800 128.600 62.600 129.000 ;
        RECT 55.800 122.800 56.400 123.000 ;
        RECT 58.800 123.000 59.600 128.600 ;
        RECT 62.000 128.200 62.600 128.600 ;
        RECT 63.800 128.800 67.400 129.400 ;
        RECT 63.800 128.200 64.400 128.800 ;
        RECT 58.800 122.800 59.400 123.000 ;
        RECT 55.800 122.200 59.400 122.800 ;
        RECT 60.400 122.800 61.200 128.000 ;
        RECT 62.000 123.400 62.800 128.200 ;
        RECT 63.600 122.800 64.400 128.200 ;
        RECT 60.400 122.200 64.400 122.800 ;
        RECT 66.800 128.200 67.400 128.800 ;
        RECT 66.800 122.200 67.600 128.200 ;
        RECT 70.000 122.200 70.800 135.700 ;
        RECT 71.600 135.600 72.400 135.700 ;
        RECT 73.400 132.400 74.000 135.800 ;
        RECT 78.200 135.400 81.800 135.800 ;
        RECT 78.800 134.400 79.600 134.800 ;
        RECT 83.000 134.400 83.600 135.800 ;
        RECT 74.800 132.800 75.600 134.400 ;
        RECT 78.000 133.800 79.600 134.400 ;
        RECT 81.200 133.800 83.600 134.400 ;
        RECT 78.000 133.600 78.800 133.800 ;
        RECT 81.200 133.600 82.000 133.800 ;
        RECT 71.600 132.200 72.400 132.400 ;
        RECT 73.200 132.200 74.000 132.400 ;
        RECT 76.400 132.200 77.200 132.400 ;
        RECT 71.600 131.600 74.000 132.200 ;
        RECT 75.600 131.600 77.200 132.200 ;
        RECT 79.600 131.600 80.400 133.200 ;
        RECT 71.800 130.200 72.400 131.600 ;
        RECT 75.600 131.200 76.400 131.600 ;
        RECT 81.200 130.200 81.800 133.600 ;
        RECT 82.800 131.600 83.600 133.200 ;
        RECT 84.400 132.800 85.200 134.400 ;
        RECT 87.600 132.800 88.400 134.400 ;
        RECT 89.200 134.300 89.800 135.800 ;
        RECT 90.800 135.700 93.200 136.300 ;
        RECT 90.800 135.600 91.600 135.700 ;
        RECT 90.800 134.300 91.600 134.400 ;
        RECT 89.200 133.700 91.600 134.300 ;
        RECT 86.000 132.200 86.800 132.400 ;
        RECT 89.200 132.200 89.800 133.700 ;
        RECT 90.800 133.600 91.600 133.700 ;
        RECT 90.800 132.200 91.600 132.400 ;
        RECT 86.000 131.600 87.600 132.200 ;
        RECT 89.200 131.600 91.600 132.200 ;
        RECT 86.800 131.200 87.600 131.600 ;
        RECT 90.800 130.200 91.400 131.600 ;
        RECT 71.600 122.200 72.400 130.200 ;
        RECT 73.200 129.600 77.200 130.200 ;
        RECT 73.200 122.200 74.000 129.600 ;
        RECT 76.400 122.200 77.200 129.600 ;
        RECT 80.600 122.200 82.600 130.200 ;
        RECT 86.000 129.600 90.000 130.200 ;
        RECT 86.000 122.200 86.800 129.600 ;
        RECT 89.200 122.200 90.000 129.600 ;
        RECT 90.800 122.200 91.600 130.200 ;
        RECT 92.400 122.200 93.200 135.700 ;
        RECT 95.600 135.800 96.400 139.800 ;
        RECT 100.000 136.200 101.600 139.800 ;
        RECT 95.600 135.200 97.800 135.800 ;
        RECT 98.800 135.400 100.400 135.600 ;
        RECT 97.000 135.000 97.800 135.200 ;
        RECT 98.400 134.800 100.400 135.400 ;
        RECT 98.400 134.400 99.000 134.800 ;
        RECT 95.600 133.800 99.000 134.400 ;
        RECT 95.600 133.600 97.200 133.800 ;
        RECT 99.600 133.400 100.400 134.200 ;
        RECT 99.600 132.800 100.200 133.400 ;
        RECT 97.600 132.200 100.200 132.800 ;
        RECT 101.000 132.800 101.600 136.200 ;
        RECT 105.200 135.800 106.000 139.800 ;
        RECT 102.200 134.800 103.000 135.600 ;
        RECT 103.600 135.200 106.000 135.800 ;
        RECT 108.400 137.800 109.200 139.800 ;
        RECT 103.600 135.000 104.400 135.200 ;
        RECT 102.400 134.400 103.000 134.800 ;
        RECT 108.400 134.400 109.000 137.800 ;
        RECT 102.400 133.600 103.200 134.400 ;
        RECT 108.400 133.600 109.200 134.400 ;
        RECT 101.000 132.400 102.000 132.800 ;
        RECT 101.000 132.200 102.800 132.400 ;
        RECT 97.600 132.000 98.400 132.200 ;
        RECT 101.400 131.600 102.800 132.200 ;
        RECT 108.400 132.300 109.000 133.600 ;
        RECT 110.000 132.300 110.800 132.400 ;
        RECT 108.400 131.700 110.800 132.300 ;
        RECT 99.800 131.400 100.600 131.600 ;
        RECT 97.200 130.800 100.600 131.400 ;
        RECT 97.200 130.200 97.800 130.800 ;
        RECT 101.400 130.200 102.000 131.600 ;
        RECT 108.400 130.200 109.000 131.700 ;
        RECT 110.000 131.600 110.800 131.700 ;
        RECT 95.600 129.600 97.800 130.200 ;
        RECT 95.600 122.200 96.400 129.600 ;
        RECT 97.000 129.400 97.800 129.600 ;
        RECT 100.000 129.600 102.000 130.200 ;
        RECT 103.600 129.600 106.000 130.200 ;
        RECT 100.000 122.200 101.600 129.600 ;
        RECT 103.600 129.400 104.400 129.600 ;
        RECT 105.200 122.200 106.000 129.600 ;
        RECT 107.400 129.400 109.200 130.200 ;
        RECT 107.400 122.200 108.200 129.400 ;
        RECT 111.600 122.200 112.400 139.800 ;
        RECT 119.600 137.800 120.400 139.800 ;
        RECT 122.800 138.400 123.600 139.800 ;
        RECT 119.200 137.600 120.400 137.800 ;
        RECT 122.600 137.800 123.600 138.400 ;
        RECT 122.600 137.600 123.200 137.800 ;
        RECT 119.200 137.000 123.200 137.600 ;
        RECT 119.200 134.400 119.800 137.000 ;
        RECT 123.400 135.600 125.200 136.400 ;
        RECT 132.400 135.200 133.200 139.800 ;
        RECT 137.200 135.200 138.000 139.800 ;
        RECT 142.000 135.200 142.800 139.800 ;
        RECT 146.800 135.200 147.600 139.800 ;
        RECT 151.600 135.200 152.400 139.800 ;
        RECT 156.400 135.200 157.200 139.800 ;
        RECT 161.200 135.200 162.000 139.800 ;
        RECT 166.000 135.200 166.800 139.800 ;
        RECT 170.800 135.200 171.600 139.800 ;
        RECT 177.200 137.800 178.000 139.800 ;
        RECT 132.400 134.600 134.600 135.200 ;
        RECT 137.200 134.600 139.400 135.200 ;
        RECT 142.000 134.600 144.200 135.200 ;
        RECT 146.800 134.600 149.000 135.200 ;
        RECT 151.600 134.600 153.800 135.200 ;
        RECT 156.400 134.600 158.600 135.200 ;
        RECT 161.200 134.600 163.400 135.200 ;
        RECT 166.000 134.600 168.200 135.200 ;
        RECT 170.800 134.600 173.000 135.200 ;
        RECT 119.200 133.600 120.400 134.400 ;
        RECT 122.000 133.600 123.600 134.400 ;
        RECT 119.200 130.400 119.800 133.600 ;
        RECT 120.400 131.600 122.000 132.400 ;
        RECT 127.600 132.300 128.400 132.400 ;
        RECT 132.400 132.300 133.200 133.200 ;
        RECT 127.600 131.700 133.200 132.300 ;
        RECT 127.600 131.600 128.400 131.700 ;
        RECT 132.400 131.600 133.200 131.700 ;
        RECT 134.000 131.600 134.600 134.600 ;
        RECT 137.200 131.600 138.000 133.200 ;
        RECT 138.800 131.600 139.400 134.600 ;
        RECT 143.600 131.600 144.200 134.600 ;
        RECT 146.800 131.600 147.600 133.200 ;
        RECT 148.400 131.600 149.000 134.600 ;
        RECT 153.200 131.600 153.800 134.600 ;
        RECT 158.000 131.600 158.600 134.600 ;
        RECT 162.800 131.600 163.400 134.600 ;
        RECT 167.600 131.600 168.200 134.600 ;
        RECT 172.400 131.600 173.000 134.600 ;
        RECT 177.200 134.400 177.800 137.800 ;
        RECT 177.200 133.600 178.000 134.400 ;
        RECT 116.400 129.800 119.800 130.400 ;
        RECT 134.000 130.800 135.200 131.600 ;
        RECT 138.800 130.800 140.000 131.600 ;
        RECT 143.600 130.800 144.800 131.600 ;
        RECT 148.400 130.800 149.600 131.600 ;
        RECT 153.200 130.800 154.400 131.600 ;
        RECT 158.000 130.800 159.200 131.600 ;
        RECT 162.800 130.800 164.000 131.600 ;
        RECT 167.600 130.800 168.800 131.600 ;
        RECT 172.400 130.800 173.600 131.600 ;
        RECT 134.000 130.200 134.600 130.800 ;
        RECT 138.800 130.200 139.400 130.800 ;
        RECT 143.600 130.200 144.200 130.800 ;
        RECT 148.400 130.200 149.000 130.800 ;
        RECT 153.200 130.200 153.800 130.800 ;
        RECT 158.000 130.200 158.600 130.800 ;
        RECT 162.800 130.200 163.400 130.800 ;
        RECT 167.600 130.200 168.200 130.800 ;
        RECT 172.400 130.200 173.000 130.800 ;
        RECT 177.200 130.200 177.800 133.600 ;
        RECT 116.400 129.600 117.200 129.800 ;
        RECT 116.600 129.000 117.200 129.600 ;
        RECT 132.400 129.600 134.600 130.200 ;
        RECT 137.200 129.600 139.400 130.200 ;
        RECT 142.000 129.600 144.200 130.200 ;
        RECT 146.800 129.600 149.000 130.200 ;
        RECT 151.600 129.600 153.800 130.200 ;
        RECT 156.400 129.600 158.600 130.200 ;
        RECT 161.200 129.600 163.400 130.200 ;
        RECT 166.000 129.600 168.200 130.200 ;
        RECT 170.800 129.600 173.000 130.200 ;
        RECT 118.200 129.000 121.800 129.200 ;
        RECT 114.800 123.000 115.600 129.000 ;
        RECT 116.400 123.400 117.200 129.000 ;
        RECT 118.000 128.600 121.800 129.000 ;
        RECT 115.000 122.800 115.600 123.000 ;
        RECT 118.000 123.000 118.800 128.600 ;
        RECT 121.200 128.200 121.800 128.600 ;
        RECT 123.000 128.800 126.600 129.400 ;
        RECT 123.000 128.200 123.600 128.800 ;
        RECT 118.000 122.800 118.600 123.000 ;
        RECT 115.000 122.200 118.600 122.800 ;
        RECT 119.600 122.800 120.400 128.000 ;
        RECT 121.200 123.400 122.000 128.200 ;
        RECT 122.800 122.800 123.600 128.200 ;
        RECT 119.600 122.200 123.600 122.800 ;
        RECT 126.000 128.200 126.600 128.800 ;
        RECT 126.000 122.200 126.800 128.200 ;
        RECT 132.400 122.200 133.200 129.600 ;
        RECT 137.200 122.200 138.000 129.600 ;
        RECT 142.000 122.200 142.800 129.600 ;
        RECT 146.800 122.200 147.600 129.600 ;
        RECT 151.600 122.200 152.400 129.600 ;
        RECT 156.400 122.200 157.200 129.600 ;
        RECT 161.200 122.200 162.000 129.600 ;
        RECT 166.000 122.200 166.800 129.600 ;
        RECT 170.800 122.200 171.600 129.600 ;
        RECT 176.200 129.400 178.000 130.200 ;
        RECT 176.200 124.400 177.000 129.400 ;
        RECT 175.600 123.600 177.000 124.400 ;
        RECT 176.200 122.200 177.000 123.600 ;
        RECT 1.200 106.800 2.000 108.400 ;
        RECT 2.800 106.200 3.600 119.800 ;
        RECT 6.600 114.400 7.400 119.800 ;
        RECT 6.000 113.600 7.400 114.400 ;
        RECT 4.400 111.600 5.200 113.200 ;
        RECT 6.600 112.600 7.400 113.600 ;
        RECT 6.600 111.800 8.400 112.600 ;
        RECT 7.600 108.400 8.200 111.800 ;
        RECT 7.600 107.600 8.400 108.400 ;
        RECT 2.800 105.600 4.600 106.200 ;
        RECT 3.800 104.400 4.600 105.600 ;
        RECT 3.800 103.600 5.200 104.400 ;
        RECT 7.600 104.200 8.200 107.600 ;
        RECT 10.800 104.800 11.600 106.400 ;
        RECT 3.800 102.200 4.600 103.600 ;
        RECT 7.600 102.200 8.400 104.200 ;
        RECT 12.400 102.200 13.200 119.800 ;
        RECT 16.200 112.400 17.000 119.800 ;
        RECT 22.000 115.800 22.800 119.800 ;
        RECT 16.000 111.800 17.000 112.400 ;
        RECT 16.000 108.400 16.600 111.800 ;
        RECT 22.200 111.600 22.800 115.800 ;
        RECT 25.200 111.800 26.000 119.800 ;
        RECT 26.800 112.400 27.600 119.800 ;
        RECT 28.400 112.400 29.200 112.600 ;
        RECT 31.200 112.400 32.800 119.800 ;
        RECT 26.800 111.800 29.200 112.400 ;
        RECT 30.800 111.800 32.800 112.400 ;
        RECT 35.000 112.400 35.800 112.600 ;
        RECT 36.400 112.400 37.200 119.800 ;
        RECT 35.000 111.800 37.200 112.400 ;
        RECT 38.000 112.400 38.800 119.800 ;
        RECT 41.200 119.200 45.200 119.800 ;
        RECT 41.200 112.400 42.000 119.200 ;
        RECT 38.000 111.800 42.000 112.400 ;
        RECT 42.800 111.800 43.600 118.600 ;
        RECT 44.400 111.800 45.200 119.200 ;
        RECT 50.800 112.400 51.600 119.800 ;
        RECT 54.000 112.400 54.800 119.800 ;
        RECT 50.800 111.800 54.800 112.400 ;
        RECT 55.600 111.800 56.400 119.800 ;
        RECT 22.200 111.000 24.600 111.600 ;
        RECT 17.200 108.800 18.000 110.400 ;
        RECT 22.000 109.600 22.800 110.400 ;
        RECT 14.000 107.600 16.600 108.400 ;
        RECT 18.800 108.200 19.600 108.400 ;
        RECT 18.000 107.600 19.600 108.200 ;
        RECT 20.400 107.600 21.200 109.200 ;
        RECT 22.200 108.800 22.800 109.600 ;
        RECT 22.200 108.200 23.200 108.800 ;
        RECT 22.400 108.000 23.200 108.200 ;
        RECT 24.000 107.600 24.600 111.000 ;
        RECT 25.400 110.400 26.000 111.800 ;
        RECT 30.800 110.400 31.400 111.800 ;
        RECT 35.000 111.200 35.600 111.800 ;
        RECT 42.800 111.200 43.400 111.800 ;
        RECT 32.200 110.600 35.600 111.200 ;
        RECT 32.200 110.400 33.000 110.600 ;
        RECT 38.800 110.400 39.600 110.800 ;
        RECT 41.400 110.600 43.400 111.200 ;
        RECT 41.400 110.400 42.000 110.600 ;
        RECT 25.200 109.600 26.000 110.400 ;
        RECT 30.000 109.800 31.400 110.400 ;
        RECT 34.400 109.800 35.200 110.000 ;
        RECT 30.000 109.600 31.800 109.800 ;
        RECT 14.200 106.200 14.800 107.600 ;
        RECT 18.000 107.200 18.800 107.600 ;
        RECT 24.000 107.400 24.800 107.600 ;
        RECT 21.800 107.000 24.800 107.400 ;
        RECT 20.600 106.800 24.800 107.000 ;
        RECT 15.800 106.200 19.400 106.600 ;
        RECT 20.600 106.400 22.400 106.800 ;
        RECT 20.600 106.200 21.200 106.400 ;
        RECT 25.400 106.200 26.000 109.600 ;
        RECT 30.800 109.200 31.800 109.600 ;
        RECT 29.600 107.600 30.400 108.400 ;
        RECT 29.800 107.200 30.400 107.600 ;
        RECT 28.400 106.800 29.200 107.000 ;
        RECT 14.000 102.200 14.800 106.200 ;
        RECT 15.600 106.000 19.600 106.200 ;
        RECT 15.600 102.200 16.400 106.000 ;
        RECT 18.800 102.200 19.600 106.000 ;
        RECT 20.400 102.200 21.200 106.200 ;
        RECT 24.600 105.200 26.000 106.200 ;
        RECT 26.800 106.200 29.200 106.800 ;
        RECT 29.800 106.400 30.600 107.200 ;
        RECT 24.600 104.400 25.400 105.200 ;
        RECT 24.600 103.600 26.000 104.400 ;
        RECT 24.600 102.200 25.400 103.600 ;
        RECT 26.800 102.200 27.600 106.200 ;
        RECT 31.200 105.800 31.800 109.200 ;
        RECT 32.600 109.200 35.200 109.800 ;
        RECT 38.000 109.800 39.600 110.400 ;
        RECT 38.000 109.600 38.800 109.800 ;
        RECT 41.200 109.600 42.000 110.400 ;
        RECT 44.400 109.600 45.200 111.200 ;
        RECT 51.600 110.400 52.400 110.800 ;
        RECT 55.600 110.400 56.200 111.800 ;
        RECT 50.800 109.800 52.400 110.400 ;
        RECT 54.000 109.800 56.400 110.400 ;
        RECT 50.800 109.600 51.600 109.800 ;
        RECT 32.600 108.600 33.200 109.200 ;
        RECT 32.400 107.800 33.200 108.600 ;
        RECT 35.600 108.300 37.200 108.400 ;
        RECT 38.000 108.300 38.800 108.400 ;
        RECT 35.600 108.200 38.800 108.300 ;
        RECT 33.800 107.700 38.800 108.200 ;
        RECT 33.800 107.600 37.200 107.700 ;
        RECT 38.000 107.600 38.800 107.700 ;
        RECT 39.600 107.600 40.400 109.200 ;
        RECT 33.800 107.200 34.400 107.600 ;
        RECT 32.400 106.600 34.400 107.200 ;
        RECT 35.000 106.800 35.800 107.000 ;
        RECT 32.400 106.400 34.000 106.600 ;
        RECT 35.000 106.200 37.200 106.800 ;
        RECT 41.400 106.400 42.000 109.600 ;
        RECT 42.600 108.800 43.400 109.600 ;
        RECT 42.800 108.400 43.400 108.800 ;
        RECT 42.800 107.600 43.600 108.400 ;
        RECT 52.400 107.600 53.200 109.200 ;
        RECT 41.400 106.200 43.600 106.400 ;
        RECT 31.200 104.400 32.800 105.800 ;
        RECT 31.200 103.600 34.000 104.400 ;
        RECT 31.200 102.200 32.800 103.600 ;
        RECT 36.400 102.200 37.200 106.200 ;
        RECT 41.000 105.600 43.600 106.200 ;
        RECT 54.000 106.200 54.600 109.800 ;
        RECT 55.600 109.600 56.400 109.800 ;
        RECT 57.200 106.800 58.000 108.400 ;
        RECT 41.000 102.200 42.600 105.600 ;
        RECT 54.000 102.200 54.800 106.200 ;
        RECT 55.600 105.600 56.400 106.400 ;
        RECT 58.800 106.200 59.600 119.800 ;
        RECT 62.800 113.600 63.600 114.400 ;
        RECT 60.400 111.600 61.200 113.200 ;
        RECT 62.800 112.400 63.400 113.600 ;
        RECT 64.200 112.400 65.000 119.800 ;
        RECT 62.000 111.800 63.400 112.400 ;
        RECT 64.000 111.800 65.000 112.400 ;
        RECT 62.000 111.600 62.800 111.800 ;
        RECT 60.400 110.300 61.200 110.400 ;
        RECT 64.000 110.300 64.600 111.800 ;
        RECT 68.400 111.600 69.200 113.200 ;
        RECT 60.400 109.700 64.600 110.300 ;
        RECT 60.400 109.600 61.200 109.700 ;
        RECT 64.000 108.400 64.600 109.700 ;
        RECT 65.200 108.800 66.000 110.400 ;
        RECT 62.000 107.600 64.600 108.400 ;
        RECT 66.800 108.200 67.600 108.400 ;
        RECT 66.000 107.600 67.600 108.200 ;
        RECT 62.200 106.200 62.800 107.600 ;
        RECT 66.000 107.200 66.800 107.600 ;
        RECT 63.800 106.200 67.400 106.600 ;
        RECT 70.000 106.200 70.800 119.800 ;
        RECT 73.200 111.800 74.000 119.800 ;
        RECT 76.400 115.800 77.200 119.800 ;
        RECT 73.200 110.400 73.800 111.800 ;
        RECT 76.400 111.600 77.000 115.800 ;
        RECT 82.200 112.600 83.000 119.800 ;
        RECT 81.200 111.800 83.000 112.600 ;
        RECT 74.600 111.000 77.000 111.600 ;
        RECT 73.200 109.600 74.000 110.400 ;
        RECT 71.600 106.800 72.400 108.400 ;
        RECT 58.800 105.600 60.600 106.200 ;
        RECT 55.400 104.800 56.200 105.600 ;
        RECT 59.800 102.200 60.600 105.600 ;
        RECT 62.000 102.200 62.800 106.200 ;
        RECT 63.600 106.000 67.600 106.200 ;
        RECT 63.600 102.200 64.400 106.000 ;
        RECT 66.800 102.200 67.600 106.000 ;
        RECT 69.000 105.600 70.800 106.200 ;
        RECT 73.200 106.200 73.800 109.600 ;
        RECT 74.600 107.600 75.200 111.000 ;
        RECT 76.400 109.600 77.200 110.400 ;
        RECT 79.600 110.300 80.400 110.400 ;
        RECT 81.400 110.300 82.000 111.800 ;
        RECT 79.600 109.700 82.000 110.300 ;
        RECT 79.600 109.600 80.400 109.700 ;
        RECT 76.400 108.800 77.000 109.600 ;
        RECT 76.000 108.200 77.000 108.800 ;
        RECT 76.000 108.000 76.800 108.200 ;
        RECT 78.000 107.600 78.800 109.200 ;
        RECT 81.400 108.400 82.000 109.700 ;
        RECT 81.200 107.600 82.000 108.400 ;
        RECT 84.400 108.300 85.200 108.400 ;
        RECT 86.000 108.300 86.800 119.800 ;
        RECT 91.800 112.600 92.600 119.800 ;
        RECT 96.600 118.400 97.400 119.800 ;
        RECT 95.600 117.600 97.400 118.400 ;
        RECT 90.800 111.800 92.600 112.600 ;
        RECT 96.600 112.400 97.400 117.600 ;
        RECT 98.000 113.600 98.800 114.400 ;
        RECT 98.200 112.400 98.800 113.600 ;
        RECT 100.400 112.400 101.200 119.800 ;
        RECT 101.800 112.400 102.600 112.600 ;
        RECT 96.600 111.800 97.600 112.400 ;
        RECT 98.200 111.800 99.600 112.400 ;
        RECT 100.400 111.800 102.600 112.400 ;
        RECT 104.800 112.400 106.400 119.800 ;
        RECT 108.400 112.400 109.200 112.600 ;
        RECT 110.000 112.400 110.800 119.800 ;
        RECT 111.800 119.200 115.400 119.800 ;
        RECT 111.800 119.000 112.400 119.200 ;
        RECT 111.600 113.000 112.400 119.000 ;
        RECT 114.800 119.000 115.400 119.200 ;
        RECT 116.400 119.200 120.400 119.800 ;
        RECT 113.200 113.000 114.000 118.600 ;
        RECT 114.800 113.400 115.600 119.000 ;
        RECT 116.400 114.000 117.200 119.200 ;
        RECT 118.000 113.800 118.800 118.600 ;
        RECT 119.600 113.800 120.400 119.200 ;
        RECT 118.000 113.400 118.600 113.800 ;
        RECT 114.800 113.000 118.600 113.400 ;
        RECT 113.400 112.400 114.000 113.000 ;
        RECT 115.000 112.800 118.600 113.000 ;
        RECT 119.800 113.200 120.400 113.800 ;
        RECT 122.800 113.800 123.600 119.800 ;
        RECT 129.400 119.200 133.000 119.800 ;
        RECT 129.400 119.000 130.000 119.200 ;
        RECT 122.800 113.200 123.400 113.800 ;
        RECT 119.800 112.600 123.400 113.200 ;
        RECT 129.200 113.000 130.000 119.000 ;
        RECT 132.400 119.000 133.000 119.200 ;
        RECT 134.000 119.200 138.000 119.800 ;
        RECT 130.800 113.000 131.600 118.600 ;
        RECT 132.400 113.400 133.200 119.000 ;
        RECT 134.000 114.000 134.800 119.200 ;
        RECT 135.600 113.800 136.400 118.600 ;
        RECT 137.200 113.800 138.000 119.200 ;
        RECT 135.600 113.400 136.200 113.800 ;
        RECT 132.400 113.000 136.200 113.400 ;
        RECT 131.000 112.400 131.600 113.000 ;
        RECT 132.600 112.800 136.200 113.000 ;
        RECT 137.400 113.200 138.000 113.800 ;
        RECT 140.400 113.800 141.200 119.800 ;
        RECT 142.200 119.200 145.800 119.800 ;
        RECT 142.200 119.000 142.800 119.200 ;
        RECT 140.400 113.200 141.000 113.800 ;
        RECT 137.400 112.600 141.000 113.200 ;
        RECT 142.000 113.000 142.800 119.000 ;
        RECT 145.200 119.000 145.800 119.200 ;
        RECT 146.800 119.200 150.800 119.800 ;
        RECT 143.600 113.000 144.400 118.600 ;
        RECT 145.200 113.400 146.000 119.000 ;
        RECT 146.800 114.000 147.600 119.200 ;
        RECT 148.400 113.800 149.200 118.600 ;
        RECT 150.000 113.800 150.800 119.200 ;
        RECT 148.400 113.400 149.000 113.800 ;
        RECT 145.200 113.000 149.000 113.400 ;
        RECT 143.800 112.400 144.400 113.000 ;
        RECT 145.400 112.800 149.000 113.000 ;
        RECT 150.200 113.200 150.800 113.800 ;
        RECT 153.200 113.800 154.000 119.800 ;
        RECT 153.200 113.200 153.800 113.800 ;
        RECT 150.200 112.600 153.800 113.200 ;
        RECT 104.800 111.800 106.800 112.400 ;
        RECT 108.400 111.800 110.800 112.400 ;
        RECT 113.200 112.200 114.000 112.400 ;
        RECT 130.800 112.200 131.600 112.400 ;
        RECT 143.600 112.200 144.400 112.400 ;
        RECT 91.000 108.400 91.600 111.800 ;
        RECT 95.600 108.800 96.400 110.400 ;
        RECT 97.000 108.400 97.600 111.800 ;
        RECT 98.800 111.600 99.600 111.800 ;
        RECT 98.900 110.300 99.500 111.600 ;
        RECT 102.000 111.200 102.600 111.800 ;
        RECT 102.000 110.600 105.400 111.200 ;
        RECT 104.600 110.400 105.400 110.600 ;
        RECT 106.200 110.400 106.800 111.800 ;
        RECT 113.200 111.600 116.600 112.200 ;
        RECT 130.800 111.600 134.200 112.200 ;
        RECT 143.600 111.600 147.000 112.200 ;
        RECT 154.800 111.600 155.600 113.200 ;
        RECT 106.200 110.300 107.600 110.400 ;
        RECT 113.200 110.300 114.000 110.400 ;
        RECT 98.900 109.700 101.100 110.300 ;
        RECT 100.500 108.400 101.100 109.700 ;
        RECT 102.400 109.800 103.200 110.000 ;
        RECT 106.200 109.800 114.000 110.300 ;
        RECT 102.400 109.200 105.000 109.800 ;
        RECT 104.400 108.600 105.000 109.200 ;
        RECT 105.800 109.700 114.000 109.800 ;
        RECT 105.800 109.600 107.600 109.700 ;
        RECT 113.200 109.600 114.000 109.700 ;
        RECT 105.800 109.200 106.800 109.600 ;
        RECT 84.400 107.700 86.800 108.300 ;
        RECT 84.400 107.600 85.200 107.700 ;
        RECT 74.400 107.400 75.200 107.600 ;
        RECT 74.400 107.000 77.400 107.400 ;
        RECT 74.400 106.800 78.600 107.000 ;
        RECT 76.800 106.400 78.600 106.800 ;
        RECT 78.000 106.200 78.600 106.400 ;
        RECT 69.000 102.200 69.800 105.600 ;
        RECT 73.200 105.200 74.600 106.200 ;
        RECT 73.800 104.400 74.600 105.200 ;
        RECT 73.200 103.600 74.600 104.400 ;
        RECT 73.800 102.200 74.600 103.600 ;
        RECT 78.000 102.200 78.800 106.200 ;
        RECT 79.600 104.800 80.400 106.400 ;
        RECT 81.400 104.200 82.000 107.600 ;
        RECT 86.000 106.200 86.800 107.700 ;
        RECT 90.800 107.600 91.600 108.400 ;
        RECT 92.400 108.300 93.200 108.400 ;
        RECT 94.000 108.300 94.800 108.400 ;
        RECT 92.400 108.200 94.800 108.300 ;
        RECT 92.400 107.700 95.600 108.200 ;
        RECT 92.400 107.600 93.200 107.700 ;
        RECT 94.000 107.600 95.600 107.700 ;
        RECT 97.000 107.600 99.600 108.400 ;
        RECT 100.400 108.200 102.000 108.400 ;
        RECT 100.400 107.600 103.800 108.200 ;
        RECT 104.400 107.800 105.200 108.600 ;
        RECT 91.000 106.400 91.600 107.600 ;
        RECT 94.800 107.200 95.600 107.600 ;
        RECT 81.200 102.200 82.000 104.200 ;
        RECT 85.000 105.600 86.800 106.200 ;
        RECT 90.800 105.600 91.600 106.400 ;
        RECT 94.200 106.200 97.800 106.600 ;
        RECT 98.800 106.200 99.400 107.600 ;
        RECT 103.200 107.200 103.800 107.600 ;
        RECT 101.800 106.800 102.600 107.000 ;
        RECT 100.400 106.200 102.600 106.800 ;
        RECT 103.200 106.600 105.200 107.200 ;
        RECT 103.600 106.400 105.200 106.600 ;
        RECT 85.000 102.200 85.800 105.600 ;
        RECT 91.000 104.200 91.600 105.600 ;
        RECT 90.800 102.200 91.600 104.200 ;
        RECT 94.000 106.000 98.000 106.200 ;
        RECT 94.000 102.200 94.800 106.000 ;
        RECT 97.200 102.200 98.000 106.000 ;
        RECT 98.800 102.200 99.600 106.200 ;
        RECT 100.400 102.200 101.200 106.200 ;
        RECT 105.800 105.800 106.400 109.200 ;
        RECT 107.200 107.600 108.000 108.400 ;
        RECT 109.200 108.300 110.800 108.400 ;
        RECT 111.600 108.300 112.400 108.400 ;
        RECT 109.200 107.700 112.400 108.300 ;
        RECT 109.200 107.600 110.800 107.700 ;
        RECT 111.600 107.600 112.400 107.700 ;
        RECT 107.200 107.200 107.800 107.600 ;
        RECT 107.000 106.400 107.800 107.200 ;
        RECT 108.400 106.800 109.200 107.000 ;
        RECT 108.400 106.200 110.800 106.800 ;
        RECT 104.800 102.200 106.400 105.800 ;
        RECT 110.000 102.200 110.800 106.200 ;
        RECT 116.000 105.000 116.600 111.600 ;
        RECT 117.200 110.300 118.800 110.400 ;
        RECT 121.200 110.300 122.000 110.400 ;
        RECT 117.200 109.700 122.000 110.300 ;
        RECT 117.200 109.600 118.800 109.700 ;
        RECT 121.200 109.600 122.000 109.700 ;
        RECT 118.800 107.600 120.400 108.400 ;
        RECT 118.000 106.300 118.800 106.400 ;
        RECT 120.200 106.300 122.000 106.400 ;
        RECT 124.400 106.300 125.200 106.400 ;
        RECT 118.000 105.700 125.200 106.300 ;
        RECT 118.000 105.600 118.800 105.700 ;
        RECT 120.200 105.600 122.000 105.700 ;
        RECT 124.400 105.600 125.200 105.700 ;
        RECT 133.600 105.000 134.200 111.600 ;
        RECT 145.200 111.400 147.000 111.600 ;
        RECT 134.800 109.600 136.400 110.400 ;
        RECT 136.400 107.600 138.000 108.400 ;
        RECT 135.600 106.300 136.400 106.400 ;
        RECT 137.800 106.300 139.600 106.400 ;
        RECT 135.600 105.700 139.600 106.300 ;
        RECT 135.600 105.600 136.400 105.700 ;
        RECT 137.800 105.600 139.600 105.700 ;
        RECT 146.400 105.000 147.000 111.400 ;
        RECT 147.600 109.600 149.200 110.400 ;
        RECT 149.200 107.600 150.800 108.400 ;
        RECT 148.400 106.300 149.200 106.400 ;
        RECT 150.600 106.300 152.400 106.400 ;
        RECT 148.400 105.700 152.400 106.300 ;
        RECT 156.400 106.200 157.200 119.800 ;
        RECT 159.600 111.800 160.400 119.800 ;
        RECT 162.800 115.800 163.600 119.800 ;
        RECT 159.600 110.400 160.200 111.800 ;
        RECT 162.800 111.600 163.400 115.800 ;
        RECT 166.000 112.400 166.800 119.800 ;
        RECT 173.400 112.600 174.200 119.800 ;
        RECT 166.000 111.800 168.200 112.400 ;
        RECT 172.400 111.800 174.200 112.600 ;
        RECT 161.000 111.000 163.400 111.600 ;
        RECT 167.600 111.200 168.200 111.800 ;
        RECT 159.600 109.600 160.400 110.400 ;
        RECT 158.000 106.800 158.800 108.400 ;
        RECT 148.400 105.600 149.200 105.700 ;
        RECT 150.600 105.600 152.400 105.700 ;
        RECT 155.400 105.600 157.200 106.200 ;
        RECT 159.600 106.200 160.200 109.600 ;
        RECT 161.000 107.600 161.600 111.000 ;
        RECT 167.600 110.400 168.800 111.200 ;
        RECT 162.800 109.600 163.600 110.400 ;
        RECT 162.800 108.800 163.400 109.600 ;
        RECT 162.400 108.200 163.400 108.800 ;
        RECT 162.400 108.000 163.200 108.200 ;
        RECT 164.400 107.600 165.200 109.200 ;
        RECT 166.000 108.800 166.800 110.400 ;
        RECT 160.800 107.400 161.600 107.600 ;
        RECT 167.600 107.400 168.200 110.400 ;
        RECT 172.600 108.400 173.200 111.800 ;
        RECT 170.800 108.300 171.600 108.400 ;
        RECT 172.400 108.300 173.200 108.400 ;
        RECT 170.800 107.700 173.200 108.300 ;
        RECT 170.800 107.600 171.600 107.700 ;
        RECT 172.400 107.600 173.200 107.700 ;
        RECT 160.800 107.000 163.800 107.400 ;
        RECT 160.800 106.800 165.000 107.000 ;
        RECT 163.200 106.400 165.000 106.800 ;
        RECT 164.400 106.200 165.000 106.400 ;
        RECT 166.000 106.800 168.200 107.400 ;
        RECT 116.000 104.400 120.000 105.000 ;
        RECT 116.000 104.200 117.200 104.400 ;
        RECT 116.400 102.200 117.200 104.200 ;
        RECT 119.400 104.200 120.000 104.400 ;
        RECT 133.600 104.400 137.600 105.000 ;
        RECT 133.600 104.200 134.800 104.400 ;
        RECT 119.400 103.600 120.400 104.200 ;
        RECT 119.600 102.200 120.400 103.600 ;
        RECT 134.000 102.200 134.800 104.200 ;
        RECT 137.000 104.200 137.600 104.400 ;
        RECT 146.400 104.400 150.400 105.000 ;
        RECT 155.400 104.400 156.200 105.600 ;
        RECT 159.600 105.200 161.000 106.200 ;
        RECT 160.200 104.400 161.000 105.200 ;
        RECT 146.400 104.200 147.600 104.400 ;
        RECT 137.000 103.600 138.000 104.200 ;
        RECT 137.200 102.200 138.000 103.600 ;
        RECT 146.800 102.200 147.600 104.200 ;
        RECT 149.800 104.200 150.400 104.400 ;
        RECT 149.800 103.600 150.800 104.200 ;
        RECT 154.800 103.600 156.200 104.400 ;
        RECT 159.600 103.600 161.000 104.400 ;
        RECT 150.000 102.200 150.800 103.600 ;
        RECT 155.400 102.200 156.200 103.600 ;
        RECT 160.200 102.200 161.000 103.600 ;
        RECT 164.400 102.200 165.200 106.200 ;
        RECT 166.000 102.200 166.800 106.800 ;
        RECT 172.600 104.200 173.200 107.600 ;
        RECT 172.400 102.200 173.200 104.200 ;
        RECT 2.800 97.600 3.600 99.800 ;
        RECT 3.000 94.400 3.600 97.600 ;
        RECT 6.000 95.800 6.800 99.800 ;
        RECT 10.200 96.800 11.000 99.800 ;
        RECT 10.200 95.800 11.600 96.800 ;
        RECT 16.200 96.000 17.000 99.000 ;
        RECT 20.400 97.000 21.200 99.000 ;
        RECT 6.200 95.600 6.800 95.800 ;
        RECT 6.200 95.200 8.000 95.600 ;
        RECT 6.200 95.000 10.400 95.200 ;
        RECT 7.400 94.600 10.400 95.000 ;
        RECT 2.800 93.600 3.600 94.400 ;
        RECT 3.000 90.200 3.600 93.600 ;
        RECT 9.600 94.400 10.400 94.600 ;
        RECT 9.600 91.000 10.200 94.400 ;
        RECT 11.000 92.400 11.600 95.800 ;
        RECT 15.400 95.400 17.000 96.000 ;
        RECT 15.400 95.000 16.200 95.400 ;
        RECT 15.400 94.400 16.000 95.000 ;
        RECT 20.600 94.800 21.200 97.000 ;
        RECT 22.000 96.000 22.800 99.800 ;
        RECT 25.200 96.000 26.000 99.800 ;
        RECT 22.000 95.800 26.000 96.000 ;
        RECT 26.800 95.800 27.600 99.800 ;
        RECT 28.400 95.800 29.200 99.800 ;
        RECT 32.800 96.200 34.400 99.800 ;
        RECT 22.200 95.400 25.800 95.800 ;
        RECT 14.000 93.600 16.000 94.400 ;
        RECT 17.000 94.200 21.200 94.800 ;
        RECT 22.800 94.400 23.600 94.800 ;
        RECT 26.800 94.400 27.400 95.800 ;
        RECT 28.400 95.200 30.600 95.800 ;
        RECT 31.600 95.400 33.200 95.600 ;
        RECT 29.800 95.000 30.600 95.200 ;
        RECT 31.200 94.800 33.200 95.400 ;
        RECT 31.200 94.400 31.800 94.800 ;
        RECT 17.000 93.800 18.000 94.200 ;
        RECT 10.800 92.300 11.600 92.400 ;
        RECT 14.000 92.300 14.800 92.400 ;
        RECT 10.800 91.700 14.800 92.300 ;
        RECT 10.800 91.600 11.600 91.700 ;
        RECT 7.800 90.400 10.200 91.000 ;
        RECT 2.800 89.400 4.600 90.200 ;
        RECT 3.800 82.200 4.600 89.400 ;
        RECT 7.800 86.200 8.400 90.400 ;
        RECT 11.000 90.200 11.600 91.600 ;
        RECT 14.000 90.800 14.800 91.700 ;
        RECT 7.600 82.200 8.400 86.200 ;
        RECT 10.800 82.200 11.600 90.200 ;
        RECT 15.400 90.400 16.000 93.600 ;
        RECT 16.600 93.000 18.000 93.800 ;
        RECT 22.000 93.800 23.600 94.400 ;
        RECT 22.000 93.600 22.800 93.800 ;
        RECT 25.000 93.600 27.600 94.400 ;
        RECT 28.400 93.800 31.800 94.400 ;
        RECT 28.400 93.600 30.000 93.800 ;
        RECT 17.400 91.000 18.000 93.000 ;
        RECT 18.800 91.600 19.600 93.200 ;
        RECT 20.400 91.600 21.200 93.200 ;
        RECT 23.600 91.600 24.400 93.200 ;
        RECT 25.000 92.300 25.600 93.600 ;
        RECT 32.400 93.400 33.200 94.200 ;
        RECT 32.400 92.800 33.000 93.400 ;
        RECT 28.400 92.300 29.200 92.400 ;
        RECT 25.000 91.700 29.200 92.300 ;
        RECT 30.400 92.200 33.000 92.800 ;
        RECT 33.800 92.800 34.400 96.200 ;
        RECT 38.000 95.800 38.800 99.800 ;
        RECT 35.000 94.800 35.800 95.600 ;
        RECT 36.400 95.200 38.800 95.800 ;
        RECT 36.400 95.000 37.200 95.200 ;
        RECT 35.200 94.400 35.800 94.800 ;
        RECT 35.200 93.600 36.000 94.400 ;
        RECT 33.800 92.400 34.800 92.800 ;
        RECT 33.800 92.200 35.600 92.400 ;
        RECT 30.400 92.000 31.200 92.200 ;
        RECT 17.400 90.400 21.200 91.000 ;
        RECT 15.400 89.800 16.400 90.400 ;
        RECT 15.400 89.200 17.000 89.800 ;
        RECT 16.200 82.200 17.000 89.200 ;
        RECT 20.600 87.000 21.200 90.400 ;
        RECT 25.000 90.200 25.600 91.700 ;
        RECT 28.400 91.600 29.200 91.700 ;
        RECT 34.200 91.600 35.600 92.200 ;
        RECT 32.600 91.400 33.400 91.600 ;
        RECT 30.000 90.800 33.400 91.400 ;
        RECT 26.800 90.200 27.600 90.400 ;
        RECT 30.000 90.200 30.600 90.800 ;
        RECT 34.200 90.400 34.800 91.600 ;
        RECT 34.200 90.200 35.600 90.400 ;
        RECT 41.200 90.300 42.000 99.800 ;
        RECT 46.400 94.400 47.200 99.800 ;
        RECT 46.000 94.200 47.200 94.400 ;
        RECT 55.200 94.200 56.000 99.800 ;
        RECT 63.000 96.400 63.800 99.800 ;
        RECT 62.000 95.800 63.800 96.400 ;
        RECT 46.000 93.600 48.200 94.200 ;
        RECT 44.400 91.600 46.000 92.400 ;
        RECT 42.800 90.300 43.600 91.200 ;
        RECT 20.400 83.000 21.200 87.000 ;
        RECT 24.600 89.600 25.600 90.200 ;
        RECT 26.200 89.600 27.600 90.200 ;
        RECT 28.400 89.600 30.600 90.200 ;
        RECT 24.600 82.200 25.400 89.600 ;
        RECT 26.200 88.400 26.800 89.600 ;
        RECT 26.000 87.600 26.800 88.400 ;
        RECT 28.400 82.200 29.200 89.600 ;
        RECT 29.800 89.400 30.600 89.600 ;
        RECT 32.800 89.600 35.600 90.200 ;
        RECT 36.400 89.600 38.800 90.200 ;
        RECT 32.800 82.200 34.400 89.600 ;
        RECT 36.400 89.400 37.200 89.600 ;
        RECT 38.000 82.200 38.800 89.600 ;
        RECT 41.200 89.700 43.600 90.300 ;
        RECT 41.200 82.200 42.000 89.700 ;
        RECT 42.800 89.600 43.600 89.700 ;
        RECT 47.600 90.400 48.200 93.600 ;
        RECT 54.200 93.800 56.000 94.200 ;
        RECT 54.200 93.600 55.800 93.800 ;
        RECT 60.400 93.600 61.200 95.200 ;
        RECT 54.200 90.400 54.800 93.600 ;
        RECT 55.600 91.600 58.000 92.400 ;
        RECT 47.600 89.600 48.400 90.400 ;
        RECT 54.000 89.600 54.800 90.400 ;
        RECT 58.800 89.600 59.600 91.200 ;
        RECT 46.000 87.600 46.800 89.200 ;
        RECT 47.600 87.000 48.200 89.600 ;
        RECT 44.600 86.400 48.200 87.000 ;
        RECT 44.600 86.200 45.200 86.400 ;
        RECT 44.400 82.200 45.200 86.200 ;
        RECT 47.600 86.200 48.200 86.400 ;
        RECT 54.200 87.000 54.800 89.600 ;
        RECT 55.600 87.600 56.400 89.200 ;
        RECT 54.200 86.400 57.800 87.000 ;
        RECT 54.200 86.200 54.800 86.400 ;
        RECT 47.600 82.200 48.400 86.200 ;
        RECT 54.000 82.200 54.800 86.200 ;
        RECT 57.200 86.200 57.800 86.400 ;
        RECT 57.200 82.200 58.000 86.200 ;
        RECT 62.000 82.200 62.800 95.800 ;
        RECT 68.800 94.200 69.600 99.800 ;
        RECT 71.600 98.300 72.400 98.400 ;
        RECT 76.400 98.300 77.200 99.800 ;
        RECT 79.600 98.400 80.400 99.800 ;
        RECT 71.600 97.700 77.200 98.300 ;
        RECT 71.600 97.600 72.400 97.700 ;
        RECT 76.000 97.600 77.200 97.700 ;
        RECT 79.400 97.800 80.400 98.400 ;
        RECT 79.400 97.600 80.000 97.800 ;
        RECT 76.000 97.000 80.000 97.600 ;
        RECT 68.800 93.800 70.600 94.200 ;
        RECT 69.000 93.600 70.600 93.800 ;
        RECT 66.800 91.600 68.400 92.400 ;
        RECT 63.600 90.300 64.400 90.400 ;
        RECT 65.200 90.300 66.000 91.200 ;
        RECT 63.600 89.700 66.000 90.300 ;
        RECT 63.600 88.800 64.400 89.700 ;
        RECT 65.200 89.600 66.000 89.700 ;
        RECT 70.000 90.400 70.600 93.600 ;
        RECT 76.000 90.400 76.600 97.000 ;
        RECT 78.800 94.300 80.400 94.400 ;
        RECT 84.400 94.300 85.200 99.800 ;
        RECT 89.200 97.800 90.000 99.800 ;
        RECT 95.600 98.400 96.400 99.800 ;
        RECT 86.000 95.600 86.800 97.200 ;
        RECT 89.200 94.400 89.800 97.800 ;
        RECT 95.600 97.600 96.600 98.400 ;
        RECT 98.800 97.800 99.600 99.800 ;
        RECT 102.000 98.300 102.800 98.400 ;
        RECT 105.200 98.300 106.000 99.800 ;
        RECT 98.800 97.600 100.000 97.800 ;
        RECT 102.000 97.700 106.000 98.300 ;
        RECT 102.000 97.600 102.800 97.700 ;
        RECT 90.800 96.300 91.600 97.200 ;
        RECT 96.000 97.000 100.000 97.600 ;
        RECT 94.000 96.300 96.400 96.400 ;
        RECT 90.800 95.700 96.400 96.300 ;
        RECT 90.800 95.600 91.600 95.700 ;
        RECT 94.000 95.600 96.400 95.700 ;
        RECT 78.800 93.700 85.200 94.300 ;
        RECT 78.800 93.600 80.400 93.700 ;
        RECT 77.200 91.600 78.800 92.400 ;
        RECT 70.000 89.600 70.800 90.400 ;
        RECT 73.200 89.800 76.600 90.400 ;
        RECT 73.200 89.600 74.000 89.800 ;
        RECT 68.400 87.600 69.200 89.200 ;
        RECT 70.000 87.000 70.600 89.600 ;
        RECT 73.400 89.000 74.000 89.600 ;
        RECT 75.000 89.000 78.600 89.200 ;
        RECT 67.000 86.400 70.600 87.000 ;
        RECT 67.000 86.200 67.600 86.400 ;
        RECT 66.800 82.200 67.600 86.200 ;
        RECT 70.000 86.200 70.600 86.400 ;
        RECT 70.000 82.200 70.800 86.200 ;
        RECT 71.600 83.000 72.400 89.000 ;
        RECT 73.200 83.400 74.000 89.000 ;
        RECT 74.800 88.600 78.600 89.000 ;
        RECT 71.800 82.800 72.400 83.000 ;
        RECT 74.800 83.000 75.600 88.600 ;
        RECT 78.000 88.200 78.600 88.600 ;
        RECT 79.800 88.800 83.400 89.400 ;
        RECT 79.800 88.200 80.400 88.800 ;
        RECT 74.800 82.800 75.400 83.000 ;
        RECT 71.800 82.200 75.400 82.800 ;
        RECT 76.400 82.800 77.200 88.000 ;
        RECT 78.000 83.400 78.800 88.200 ;
        RECT 79.600 82.800 80.400 88.200 ;
        RECT 76.400 82.200 80.400 82.800 ;
        RECT 82.800 88.200 83.400 88.800 ;
        RECT 82.800 82.200 83.600 88.200 ;
        RECT 84.400 82.200 85.200 93.700 ;
        RECT 86.000 94.300 86.800 94.400 ;
        RECT 89.200 94.300 90.000 94.400 ;
        RECT 86.000 93.700 90.000 94.300 ;
        RECT 86.000 93.600 86.800 93.700 ;
        RECT 89.200 93.600 90.000 93.700 ;
        RECT 90.800 94.300 91.600 94.400 ;
        RECT 95.600 94.300 97.200 94.400 ;
        RECT 90.800 93.700 97.200 94.300 ;
        RECT 90.800 93.600 91.600 93.700 ;
        RECT 95.600 93.600 97.200 93.700 ;
        RECT 87.600 90.800 88.400 92.400 ;
        RECT 89.200 90.200 89.800 93.600 ;
        RECT 97.200 91.600 98.800 92.400 ;
        RECT 99.400 90.400 100.000 97.000 ;
        RECT 105.200 95.800 106.000 97.700 ;
        RECT 106.800 96.000 107.600 99.800 ;
        RECT 110.000 96.000 110.800 99.800 ;
        RECT 113.200 97.800 114.000 99.800 ;
        RECT 106.800 95.800 110.800 96.000 ;
        RECT 105.400 94.400 106.000 95.800 ;
        RECT 107.000 95.400 110.600 95.800 ;
        RECT 111.600 95.600 112.400 97.200 ;
        RECT 109.200 94.400 110.000 94.800 ;
        RECT 113.400 94.400 114.000 97.800 ;
        RECT 116.400 95.200 117.200 99.800 ;
        RECT 116.400 94.600 118.600 95.200 ;
        RECT 105.200 93.600 107.800 94.400 ;
        RECT 109.200 94.300 110.800 94.400 ;
        RECT 111.600 94.300 112.400 94.400 ;
        RECT 109.200 93.800 112.400 94.300 ;
        RECT 110.000 93.700 112.400 93.800 ;
        RECT 110.000 93.600 110.800 93.700 ;
        RECT 111.600 93.600 112.400 93.700 ;
        RECT 113.200 93.600 114.000 94.400 ;
        RECT 88.200 89.400 90.000 90.200 ;
        RECT 99.400 89.800 102.800 90.400 ;
        RECT 102.000 89.600 102.800 89.800 ;
        RECT 105.200 90.200 106.000 90.400 ;
        RECT 107.200 90.200 107.800 93.600 ;
        RECT 108.400 91.600 109.200 93.200 ;
        RECT 113.400 90.200 114.000 93.600 ;
        RECT 114.800 90.800 115.600 92.400 ;
        RECT 116.400 91.600 117.200 93.200 ;
        RECT 118.000 91.600 118.600 94.600 ;
        RECT 119.600 92.400 120.400 99.800 ;
        RECT 123.800 96.400 124.600 99.800 ;
        RECT 122.800 95.800 124.600 96.400 ;
        RECT 130.800 95.800 131.600 99.800 ;
        RECT 135.200 98.400 136.800 99.800 ;
        RECT 135.200 97.600 138.000 98.400 ;
        RECT 135.200 96.200 136.800 97.600 ;
        RECT 121.200 93.600 122.000 95.200 ;
        RECT 122.800 94.300 123.600 95.800 ;
        RECT 130.800 95.200 133.400 95.800 ;
        RECT 132.600 95.000 133.400 95.200 ;
        RECT 134.000 94.800 135.600 95.600 ;
        RECT 130.800 94.300 132.400 94.400 ;
        RECT 122.800 94.200 132.400 94.300 ;
        RECT 136.200 94.200 136.800 96.200 ;
        RECT 140.400 95.800 141.200 99.800 ;
        RECT 142.000 95.800 142.800 99.800 ;
        RECT 143.600 96.000 144.400 99.800 ;
        RECT 146.800 96.000 147.600 99.800 ;
        RECT 143.600 95.800 147.600 96.000 ;
        RECT 149.000 96.400 149.800 99.800 ;
        RECT 155.800 96.400 156.600 99.800 ;
        RECT 160.600 96.400 161.400 99.800 ;
        RECT 149.000 95.800 150.800 96.400 ;
        RECT 137.400 94.800 138.200 95.600 ;
        RECT 138.800 95.200 141.200 95.800 ;
        RECT 138.800 95.000 139.600 95.200 ;
        RECT 122.800 94.000 133.000 94.200 ;
        RECT 122.800 93.700 135.200 94.000 ;
        RECT 118.000 90.800 119.200 91.600 ;
        RECT 118.000 90.200 118.600 90.800 ;
        RECT 119.800 90.200 120.400 92.400 ;
        RECT 105.200 89.600 106.600 90.200 ;
        RECT 107.200 89.600 108.200 90.200 ;
        RECT 88.200 82.200 89.000 89.400 ;
        RECT 92.600 88.800 96.200 89.400 ;
        RECT 92.600 88.200 93.200 88.800 ;
        RECT 92.400 82.200 93.200 88.200 ;
        RECT 95.600 88.200 96.200 88.800 ;
        RECT 97.400 89.000 101.000 89.200 ;
        RECT 102.000 89.000 102.600 89.600 ;
        RECT 97.400 88.600 101.200 89.000 ;
        RECT 97.400 88.200 98.000 88.600 ;
        RECT 95.600 82.800 96.400 88.200 ;
        RECT 97.200 83.400 98.000 88.200 ;
        RECT 98.800 82.800 99.600 88.000 ;
        RECT 100.400 83.000 101.200 88.600 ;
        RECT 102.000 83.400 102.800 89.000 ;
        RECT 95.600 82.200 99.600 82.800 ;
        RECT 100.600 82.800 101.200 83.000 ;
        RECT 103.600 83.000 104.400 89.000 ;
        RECT 106.000 88.400 106.600 89.600 ;
        RECT 106.000 87.600 106.800 88.400 ;
        RECT 103.600 82.800 104.200 83.000 ;
        RECT 100.600 82.200 104.200 82.800 ;
        RECT 107.400 82.200 108.200 89.600 ;
        RECT 113.200 89.400 115.000 90.200 ;
        RECT 114.200 84.400 115.000 89.400 ;
        RECT 116.400 89.600 118.600 90.200 ;
        RECT 114.200 83.600 115.600 84.400 ;
        RECT 114.200 82.200 115.000 83.600 ;
        RECT 116.400 82.200 117.200 89.600 ;
        RECT 119.600 82.200 120.400 90.200 ;
        RECT 122.800 82.200 123.600 93.700 ;
        RECT 130.800 93.600 135.200 93.700 ;
        RECT 132.400 93.400 135.200 93.600 ;
        RECT 134.400 93.200 135.200 93.400 ;
        RECT 135.800 93.600 136.800 94.200 ;
        RECT 137.600 94.400 138.200 94.800 ;
        RECT 142.200 94.400 142.800 95.800 ;
        RECT 143.800 95.400 147.400 95.800 ;
        RECT 137.600 93.600 138.400 94.400 ;
        RECT 142.000 93.600 144.600 94.400 ;
        RECT 148.400 94.300 149.200 94.400 ;
        RECT 150.000 94.300 150.800 95.800 ;
        RECT 154.800 95.800 156.600 96.400 ;
        RECT 159.600 95.800 161.400 96.400 ;
        RECT 162.800 95.800 163.600 99.800 ;
        RECT 167.200 98.400 168.800 99.800 ;
        RECT 166.000 97.600 168.800 98.400 ;
        RECT 167.200 96.200 168.800 97.600 ;
        RECT 148.400 93.700 150.800 94.300 ;
        RECT 148.400 93.600 149.200 93.700 ;
        RECT 135.800 92.400 136.400 93.600 ;
        RECT 133.000 92.200 133.800 92.400 ;
        RECT 133.000 91.600 134.600 92.200 ;
        RECT 135.600 91.600 136.400 92.400 ;
        RECT 133.800 91.400 134.600 91.600 ;
        RECT 124.400 88.800 125.200 90.400 ;
        RECT 135.800 90.200 136.400 91.600 ;
        RECT 142.000 90.200 142.800 90.400 ;
        RECT 144.000 90.200 144.600 93.600 ;
        RECT 145.200 91.600 146.000 93.200 ;
        RECT 130.800 89.600 133.400 90.200 ;
        RECT 130.800 82.200 131.600 89.600 ;
        RECT 132.600 89.400 133.400 89.600 ;
        RECT 135.200 82.200 136.800 90.200 ;
        RECT 138.800 89.600 141.200 90.200 ;
        RECT 142.000 89.600 143.400 90.200 ;
        RECT 144.000 89.600 145.000 90.200 ;
        RECT 138.800 89.400 139.600 89.600 ;
        RECT 140.400 82.200 141.200 89.600 ;
        RECT 142.800 88.400 143.400 89.600 ;
        RECT 142.800 87.600 143.600 88.400 ;
        RECT 144.200 82.200 145.000 89.600 ;
        RECT 148.400 88.800 149.200 90.400 ;
        RECT 150.000 82.200 150.800 93.700 ;
        RECT 151.600 94.300 152.400 95.200 ;
        RECT 153.200 94.300 154.000 95.200 ;
        RECT 151.600 93.700 154.000 94.300 ;
        RECT 151.600 93.600 152.400 93.700 ;
        RECT 153.200 93.600 154.000 93.700 ;
        RECT 154.800 82.200 155.600 95.800 ;
        RECT 158.000 93.600 158.800 95.200 ;
        RECT 156.400 90.300 157.200 90.400 ;
        RECT 158.000 90.300 158.800 90.400 ;
        RECT 156.400 89.700 158.800 90.300 ;
        RECT 156.400 88.800 157.200 89.700 ;
        RECT 158.000 89.600 158.800 89.700 ;
        RECT 159.600 82.200 160.400 95.800 ;
        RECT 162.800 95.200 165.400 95.800 ;
        RECT 164.600 95.000 165.400 95.200 ;
        RECT 166.000 94.800 167.600 95.600 ;
        RECT 162.800 94.200 164.400 94.400 ;
        RECT 168.200 94.200 168.800 96.200 ;
        RECT 172.400 95.800 173.200 99.800 ;
        RECT 169.400 94.800 170.200 95.600 ;
        RECT 170.800 95.200 173.200 95.800 ;
        RECT 174.000 95.200 174.800 99.800 ;
        RECT 170.800 95.000 171.600 95.200 ;
        RECT 162.800 94.000 165.000 94.200 ;
        RECT 162.800 93.600 167.200 94.000 ;
        RECT 164.400 93.400 167.200 93.600 ;
        RECT 166.400 93.200 167.200 93.400 ;
        RECT 167.800 93.600 168.800 94.200 ;
        RECT 169.600 94.400 170.200 94.800 ;
        RECT 174.000 94.600 176.200 95.200 ;
        RECT 169.600 93.600 170.400 94.400 ;
        RECT 167.800 92.400 168.400 93.600 ;
        RECT 165.000 92.200 165.800 92.400 ;
        RECT 165.000 91.600 166.600 92.200 ;
        RECT 167.600 91.600 168.400 92.400 ;
        RECT 165.800 91.400 166.600 91.600 ;
        RECT 161.200 88.800 162.000 90.400 ;
        RECT 167.800 90.200 168.400 91.600 ;
        RECT 175.600 91.600 176.200 94.600 ;
        RECT 175.600 90.800 176.800 91.600 ;
        RECT 175.600 90.200 176.200 90.800 ;
        RECT 162.800 89.600 165.400 90.200 ;
        RECT 162.800 82.200 163.600 89.600 ;
        RECT 164.600 89.400 165.400 89.600 ;
        RECT 167.200 82.200 168.800 90.200 ;
        RECT 170.800 89.600 173.200 90.200 ;
        RECT 170.800 89.400 171.600 89.600 ;
        RECT 172.400 82.200 173.200 89.600 ;
        RECT 174.000 89.600 176.200 90.200 ;
        RECT 174.000 82.200 174.800 89.600 ;
        RECT 4.400 72.400 5.200 79.800 ;
        RECT 3.000 71.800 5.200 72.400 ;
        RECT 6.600 74.400 7.400 79.800 ;
        RECT 6.600 73.600 8.400 74.400 ;
        RECT 6.600 72.600 7.400 73.600 ;
        RECT 11.400 72.600 12.200 79.800 ;
        RECT 15.600 75.800 16.400 79.800 ;
        RECT 15.800 75.600 16.400 75.800 ;
        RECT 18.800 75.800 19.600 79.800 ;
        RECT 23.600 75.800 24.400 79.800 ;
        RECT 18.800 75.600 19.400 75.800 ;
        RECT 15.800 75.000 19.400 75.600 ;
        RECT 23.800 75.600 24.400 75.800 ;
        RECT 26.800 75.800 27.600 79.800 ;
        RECT 28.400 75.800 29.200 79.800 ;
        RECT 26.800 75.600 27.400 75.800 ;
        RECT 23.800 75.000 27.400 75.600 ;
        RECT 6.600 71.800 8.400 72.600 ;
        RECT 11.400 71.800 13.200 72.600 ;
        RECT 15.800 72.400 16.400 75.000 ;
        RECT 17.200 72.800 18.000 74.400 ;
        RECT 25.200 72.800 26.000 74.400 ;
        RECT 26.800 72.400 27.400 75.000 ;
        RECT 28.600 75.600 29.200 75.800 ;
        RECT 31.600 75.600 32.400 79.800 ;
        RECT 28.600 75.000 32.200 75.600 ;
        RECT 28.600 72.400 29.200 75.000 ;
        RECT 30.000 72.800 30.800 74.400 ;
        RECT 34.800 72.400 35.600 79.800 ;
        RECT 36.400 72.400 37.200 72.600 ;
        RECT 39.200 72.400 40.800 79.800 ;
        RECT 3.000 71.200 3.600 71.800 ;
        RECT 2.400 70.400 3.600 71.200 ;
        RECT 3.000 67.400 3.600 70.400 ;
        RECT 6.000 69.600 6.800 71.200 ;
        RECT 7.600 68.400 8.200 71.800 ;
        RECT 12.400 68.400 13.000 71.800 ;
        RECT 15.600 71.600 16.400 72.400 ;
        RECT 15.800 68.400 16.400 71.600 ;
        RECT 20.400 70.800 21.200 72.400 ;
        RECT 22.000 70.800 22.800 72.400 ;
        RECT 26.800 71.600 27.600 72.400 ;
        RECT 28.400 71.600 29.200 72.400 ;
        RECT 18.000 69.600 19.600 70.400 ;
        RECT 23.600 69.600 25.200 70.400 ;
        RECT 26.800 68.400 27.400 71.600 ;
        RECT 7.600 67.600 8.400 68.400 ;
        RECT 12.400 67.600 13.200 68.400 ;
        RECT 15.800 68.200 17.400 68.400 ;
        RECT 25.800 68.200 27.400 68.400 ;
        RECT 15.800 67.800 17.600 68.200 ;
        RECT 3.000 66.800 5.200 67.400 ;
        RECT 4.400 62.200 5.200 66.800 ;
        RECT 7.600 64.200 8.200 67.600 ;
        RECT 9.200 64.800 10.000 66.400 ;
        RECT 10.800 66.300 11.600 66.400 ;
        RECT 12.400 66.300 13.000 67.600 ;
        RECT 10.800 65.700 13.100 66.300 ;
        RECT 10.800 65.600 11.600 65.700 ;
        RECT 12.400 64.200 13.000 65.700 ;
        RECT 7.600 62.200 8.400 64.200 ;
        RECT 12.400 62.200 13.200 64.200 ;
        RECT 16.800 62.200 17.600 67.800 ;
        RECT 25.600 67.800 27.400 68.200 ;
        RECT 28.600 68.400 29.200 71.600 ;
        RECT 33.200 70.800 34.000 72.400 ;
        RECT 34.800 71.800 37.200 72.400 ;
        RECT 38.800 71.800 40.800 72.400 ;
        RECT 43.000 72.400 43.800 72.600 ;
        RECT 44.400 72.400 45.200 79.800 ;
        RECT 51.600 73.600 52.400 74.400 ;
        RECT 51.600 72.400 52.200 73.600 ;
        RECT 53.000 72.400 53.800 79.800 ;
        RECT 43.000 71.800 45.200 72.400 ;
        RECT 46.000 72.300 46.800 72.400 ;
        RECT 50.800 72.300 52.200 72.400 ;
        RECT 46.000 71.800 52.200 72.300 ;
        RECT 52.800 71.800 53.800 72.400 ;
        RECT 57.200 71.800 58.000 79.800 ;
        RECT 58.800 72.400 59.600 79.800 ;
        RECT 62.000 72.400 62.800 79.800 ;
        RECT 58.800 71.800 62.800 72.400 ;
        RECT 38.800 70.400 39.400 71.800 ;
        RECT 43.000 71.200 43.600 71.800 ;
        RECT 46.000 71.700 51.600 71.800 ;
        RECT 46.000 71.600 46.800 71.700 ;
        RECT 50.800 71.600 51.600 71.700 ;
        RECT 40.200 70.600 43.600 71.200 ;
        RECT 40.200 70.400 41.000 70.600 ;
        RECT 30.800 69.600 32.400 70.400 ;
        RECT 38.000 69.800 39.400 70.400 ;
        RECT 52.800 70.300 53.400 71.800 ;
        RECT 57.400 70.400 58.000 71.800 ;
        RECT 61.200 70.400 62.000 70.800 ;
        RECT 42.400 69.800 43.200 70.000 ;
        RECT 38.000 69.600 39.800 69.800 ;
        RECT 38.800 69.200 39.800 69.600 ;
        RECT 28.600 68.200 30.200 68.400 ;
        RECT 28.600 67.800 30.400 68.200 ;
        RECT 25.600 62.200 26.400 67.800 ;
        RECT 29.600 62.200 30.400 67.800 ;
        RECT 37.600 67.600 38.400 68.400 ;
        RECT 37.800 67.200 38.400 67.600 ;
        RECT 36.400 66.800 37.200 67.000 ;
        RECT 34.800 66.200 37.200 66.800 ;
        RECT 37.800 66.400 38.600 67.200 ;
        RECT 34.800 62.200 35.600 66.200 ;
        RECT 39.200 65.800 39.800 69.200 ;
        RECT 40.600 69.200 43.200 69.800 ;
        RECT 44.500 69.700 53.400 70.300 ;
        RECT 40.600 68.600 41.200 69.200 ;
        RECT 40.400 67.800 41.200 68.600 ;
        RECT 44.500 68.400 45.100 69.700 ;
        RECT 52.800 68.400 53.400 69.700 ;
        RECT 54.000 68.800 54.800 70.400 ;
        RECT 57.200 69.800 59.600 70.400 ;
        RECT 61.200 69.800 62.800 70.400 ;
        RECT 57.200 69.600 58.000 69.800 ;
        RECT 58.800 69.600 59.600 69.800 ;
        RECT 62.000 69.600 62.800 69.800 ;
        RECT 43.600 68.200 45.200 68.400 ;
        RECT 41.800 67.600 45.200 68.200 ;
        RECT 50.800 67.600 53.400 68.400 ;
        RECT 41.800 67.200 42.400 67.600 ;
        RECT 40.400 66.600 42.400 67.200 ;
        RECT 43.000 66.800 43.800 67.000 ;
        RECT 40.400 66.400 42.000 66.600 ;
        RECT 43.000 66.200 45.200 66.800 ;
        RECT 51.000 66.200 51.600 67.600 ;
        RECT 52.600 66.200 56.200 66.600 ;
        RECT 39.200 64.400 40.800 65.800 ;
        RECT 39.200 63.600 42.000 64.400 ;
        RECT 39.200 62.200 40.800 63.600 ;
        RECT 44.400 62.200 45.200 66.200 ;
        RECT 50.800 62.200 51.600 66.200 ;
        RECT 52.400 66.000 56.400 66.200 ;
        RECT 52.400 62.200 53.200 66.000 ;
        RECT 55.600 62.200 56.400 66.000 ;
        RECT 57.200 65.600 58.000 66.400 ;
        RECT 59.000 66.200 59.600 69.600 ;
        RECT 60.400 67.600 61.200 69.200 ;
        RECT 57.400 64.800 58.200 65.600 ;
        RECT 58.800 62.200 59.600 66.200 ;
        RECT 65.200 62.200 66.000 79.800 ;
        RECT 68.400 75.800 69.200 79.800 ;
        RECT 68.600 75.600 69.200 75.800 ;
        RECT 71.600 75.800 72.400 79.800 ;
        RECT 71.600 75.600 72.200 75.800 ;
        RECT 68.600 75.000 72.200 75.600 ;
        RECT 70.000 72.800 70.800 74.400 ;
        RECT 71.600 72.400 72.200 75.000 ;
        RECT 66.800 70.800 67.600 72.400 ;
        RECT 71.600 71.600 72.400 72.400 ;
        RECT 73.200 71.600 74.000 73.200 ;
        RECT 68.400 69.600 70.000 70.400 ;
        RECT 71.600 68.400 72.200 71.600 ;
        RECT 74.800 70.300 75.600 79.800 ;
        RECT 78.000 72.400 78.800 79.800 ;
        RECT 81.200 79.200 85.200 79.800 ;
        RECT 81.200 72.400 82.000 79.200 ;
        RECT 78.000 71.800 82.000 72.400 ;
        RECT 82.800 71.800 83.600 78.600 ;
        RECT 84.400 71.800 85.200 79.200 ;
        RECT 87.600 75.800 88.400 79.800 ;
        RECT 87.800 75.600 88.400 75.800 ;
        RECT 90.800 75.800 91.600 79.800 ;
        RECT 90.800 75.600 91.400 75.800 ;
        RECT 87.800 75.000 91.400 75.600 ;
        RECT 89.200 72.800 90.000 74.400 ;
        RECT 90.800 72.400 91.400 75.000 ;
        RECT 82.800 71.200 83.400 71.800 ;
        RECT 78.800 70.400 79.600 70.800 ;
        RECT 81.400 70.600 83.400 71.200 ;
        RECT 81.400 70.400 82.000 70.600 ;
        RECT 78.000 70.300 79.600 70.400 ;
        RECT 74.800 69.800 79.600 70.300 ;
        RECT 74.800 69.700 78.800 69.800 ;
        RECT 70.600 68.300 72.200 68.400 ;
        RECT 73.200 68.300 74.000 68.400 ;
        RECT 70.600 68.200 74.000 68.300 ;
        RECT 70.400 67.700 74.000 68.200 ;
        RECT 70.400 62.200 71.200 67.700 ;
        RECT 73.200 67.600 74.000 67.700 ;
        RECT 74.800 66.200 75.600 69.700 ;
        RECT 78.000 69.600 78.800 69.700 ;
        RECT 81.200 69.600 82.000 70.400 ;
        RECT 84.400 69.600 85.200 71.200 ;
        RECT 86.000 70.800 86.800 72.400 ;
        RECT 90.800 71.600 91.600 72.400 ;
        RECT 87.600 69.600 89.200 70.400 ;
        RECT 76.400 66.800 77.200 68.400 ;
        RECT 79.600 67.600 80.400 69.200 ;
        RECT 81.400 66.200 82.000 69.600 ;
        RECT 82.600 68.800 83.400 69.600 ;
        RECT 82.800 68.400 83.400 68.800 ;
        RECT 90.800 68.400 91.400 71.600 ;
        RECT 82.800 67.600 83.600 68.400 ;
        RECT 89.800 68.200 91.400 68.400 ;
        RECT 89.600 67.800 91.400 68.200 ;
        RECT 73.800 65.600 75.600 66.200 ;
        RECT 73.800 64.400 74.600 65.600 ;
        RECT 73.200 63.600 74.600 64.400 ;
        RECT 73.800 62.200 74.600 63.600 ;
        RECT 81.000 62.200 82.600 66.200 ;
        RECT 89.600 64.400 90.400 67.800 ;
        RECT 89.200 63.600 90.400 64.400 ;
        RECT 89.600 62.200 90.400 63.600 ;
        RECT 92.400 62.200 93.200 79.800 ;
        RECT 95.600 72.400 96.400 79.800 ;
        RECT 97.200 72.400 98.000 72.600 ;
        RECT 95.600 71.800 98.000 72.400 ;
        RECT 100.000 71.800 101.600 79.800 ;
        RECT 103.400 72.400 104.200 72.600 ;
        RECT 105.200 72.400 106.000 79.800 ;
        RECT 107.600 73.600 108.400 74.400 ;
        RECT 107.600 72.400 108.200 73.600 ;
        RECT 109.000 72.400 109.800 79.800 ;
        RECT 103.400 71.800 106.000 72.400 ;
        RECT 106.800 71.800 108.200 72.400 ;
        RECT 108.800 71.800 109.800 72.400 ;
        RECT 113.200 71.800 114.000 79.800 ;
        RECT 116.400 72.400 117.200 79.800 ;
        RECT 115.000 71.800 117.200 72.400 ;
        RECT 118.000 72.400 118.800 79.800 ;
        RECT 118.000 71.800 120.200 72.400 ;
        RECT 121.200 71.800 122.000 79.800 ;
        RECT 122.800 72.400 123.600 79.800 ;
        RECT 126.000 74.300 126.800 79.800 ;
        RECT 130.800 74.300 131.600 74.400 ;
        RECT 126.000 73.700 131.600 74.300 ;
        RECT 122.800 71.800 125.000 72.400 ;
        RECT 126.000 71.800 126.800 73.700 ;
        RECT 130.800 73.600 131.600 73.700 ;
        RECT 100.400 70.400 101.000 71.800 ;
        RECT 106.800 71.600 107.600 71.800 ;
        RECT 102.200 70.400 103.000 70.600 ;
        RECT 100.400 69.600 101.200 70.400 ;
        RECT 102.200 69.800 103.800 70.400 ;
        RECT 103.000 69.600 103.800 69.800 ;
        RECT 100.400 68.400 101.000 69.600 ;
        RECT 98.400 67.600 99.200 68.400 ;
        RECT 98.600 67.200 99.200 67.600 ;
        RECT 100.000 67.800 101.000 68.400 ;
        RECT 101.600 68.600 102.400 68.800 ;
        RECT 101.600 68.400 104.400 68.600 ;
        RECT 108.800 68.400 109.400 71.800 ;
        RECT 110.000 68.800 110.800 70.400 ;
        RECT 113.200 69.600 113.800 71.800 ;
        RECT 115.000 71.200 115.600 71.800 ;
        RECT 114.400 70.400 115.600 71.200 ;
        RECT 101.600 68.300 106.000 68.400 ;
        RECT 106.800 68.300 109.400 68.400 ;
        RECT 101.600 68.000 109.400 68.300 ;
        RECT 111.600 68.200 112.400 68.400 ;
        RECT 103.800 67.800 109.400 68.000 ;
        RECT 97.200 66.800 98.000 67.000 ;
        RECT 94.000 64.800 94.800 66.400 ;
        RECT 95.600 66.200 98.000 66.800 ;
        RECT 98.600 66.400 99.400 67.200 ;
        RECT 95.600 62.200 96.400 66.200 ;
        RECT 100.000 65.800 100.600 67.800 ;
        RECT 104.400 67.700 109.400 67.800 ;
        RECT 104.400 67.600 106.000 67.700 ;
        RECT 106.800 67.600 109.400 67.700 ;
        RECT 110.800 67.600 112.400 68.200 ;
        RECT 101.200 66.400 102.800 67.200 ;
        RECT 103.400 66.800 104.200 67.000 ;
        RECT 103.400 66.200 106.000 66.800 ;
        RECT 107.000 66.200 107.600 67.600 ;
        RECT 110.800 67.200 111.600 67.600 ;
        RECT 108.600 66.200 112.200 66.600 ;
        RECT 100.000 64.400 101.600 65.800 ;
        RECT 98.800 63.600 101.600 64.400 ;
        RECT 100.000 62.200 101.600 63.600 ;
        RECT 105.200 62.200 106.000 66.200 ;
        RECT 106.800 62.200 107.600 66.200 ;
        RECT 108.400 66.000 112.400 66.200 ;
        RECT 108.400 62.200 109.200 66.000 ;
        RECT 111.600 62.200 112.400 66.000 ;
        RECT 113.200 62.200 114.000 69.600 ;
        RECT 115.000 67.400 115.600 70.400 ;
        RECT 119.600 71.200 120.200 71.800 ;
        RECT 119.600 70.400 120.800 71.200 ;
        RECT 119.600 67.400 120.200 70.400 ;
        RECT 121.400 69.600 122.000 71.800 ;
        RECT 115.000 66.800 117.200 67.400 ;
        RECT 116.400 62.200 117.200 66.800 ;
        RECT 118.000 66.800 120.200 67.400 ;
        RECT 118.000 62.200 118.800 66.800 ;
        RECT 121.200 62.200 122.000 69.600 ;
        RECT 124.400 71.200 125.000 71.800 ;
        RECT 124.400 70.400 125.600 71.200 ;
        RECT 124.400 67.400 125.000 70.400 ;
        RECT 126.200 69.600 126.800 71.800 ;
        RECT 122.800 66.800 125.000 67.400 ;
        RECT 122.800 62.200 123.600 66.800 ;
        RECT 126.000 62.200 126.800 69.600 ;
        RECT 132.400 71.800 133.200 79.800 ;
        RECT 135.600 72.400 136.400 79.800 ;
        RECT 134.200 71.800 136.400 72.400 ;
        RECT 132.400 69.600 133.000 71.800 ;
        RECT 134.200 71.200 134.800 71.800 ;
        RECT 133.600 70.400 134.800 71.200 ;
        RECT 132.400 62.200 133.200 69.600 ;
        RECT 134.200 67.400 134.800 70.400 ;
        RECT 134.200 66.800 136.400 67.400 ;
        RECT 137.200 66.800 138.000 68.400 ;
        RECT 135.600 62.200 136.400 66.800 ;
        RECT 138.800 66.200 139.600 79.800 ;
        RECT 142.800 73.600 143.600 74.400 ;
        RECT 140.400 71.600 141.200 73.200 ;
        RECT 142.800 72.400 143.400 73.600 ;
        RECT 144.200 72.400 145.000 79.800 ;
        RECT 142.000 71.800 143.400 72.400 ;
        RECT 144.000 71.800 145.000 72.400 ;
        RECT 148.400 72.400 149.200 79.800 ;
        RECT 150.200 72.400 151.000 72.600 ;
        RECT 148.400 71.800 151.000 72.400 ;
        RECT 152.800 71.800 154.400 79.800 ;
        RECT 156.400 72.400 157.200 72.600 ;
        RECT 158.000 72.400 158.800 79.800 ;
        RECT 162.200 78.400 163.000 79.800 ;
        RECT 162.200 77.600 163.600 78.400 ;
        RECT 162.200 72.600 163.000 77.600 ;
        RECT 156.400 71.800 158.800 72.400 ;
        RECT 161.200 71.800 163.000 72.600 ;
        RECT 167.600 72.400 168.400 79.800 ;
        RECT 166.200 71.800 168.400 72.400 ;
        RECT 169.200 72.400 170.000 79.800 ;
        RECT 174.000 72.400 174.800 79.800 ;
        RECT 169.200 71.800 171.400 72.400 ;
        RECT 174.000 71.800 176.200 72.400 ;
        RECT 142.000 71.600 142.800 71.800 ;
        RECT 144.000 68.400 144.600 71.800 ;
        RECT 151.400 70.400 152.200 70.600 ;
        RECT 153.400 70.400 154.000 71.800 ;
        RECT 145.200 68.800 146.000 70.400 ;
        RECT 150.600 69.800 152.200 70.400 ;
        RECT 150.600 69.600 151.400 69.800 ;
        RECT 153.200 69.600 154.000 70.400 ;
        RECT 152.000 68.600 152.800 68.800 ;
        RECT 150.000 68.400 152.800 68.600 ;
        RECT 142.000 67.600 144.600 68.400 ;
        RECT 148.400 68.000 152.800 68.400 ;
        RECT 153.400 68.400 154.000 69.600 ;
        RECT 161.400 68.400 162.000 71.800 ;
        RECT 166.200 71.200 166.800 71.800 ;
        RECT 165.600 70.400 166.800 71.200 ;
        RECT 148.400 67.800 150.600 68.000 ;
        RECT 153.400 67.800 154.400 68.400 ;
        RECT 148.400 67.600 150.000 67.800 ;
        RECT 142.200 66.200 142.800 67.600 ;
        RECT 150.200 66.800 151.000 67.000 ;
        RECT 143.800 66.200 147.400 66.600 ;
        RECT 148.400 66.200 151.000 66.800 ;
        RECT 151.600 66.400 153.200 67.200 ;
        RECT 138.800 65.600 140.600 66.200 ;
        RECT 139.800 64.400 140.600 65.600 ;
        RECT 139.800 63.600 141.200 64.400 ;
        RECT 139.800 62.200 140.600 63.600 ;
        RECT 142.000 62.200 142.800 66.200 ;
        RECT 143.600 66.000 147.600 66.200 ;
        RECT 143.600 62.200 144.400 66.000 ;
        RECT 146.800 62.200 147.600 66.000 ;
        RECT 148.400 62.200 149.200 66.200 ;
        RECT 153.800 65.800 154.400 67.800 ;
        RECT 155.200 67.600 156.000 68.400 ;
        RECT 161.200 67.600 162.000 68.400 ;
        RECT 155.200 67.200 155.800 67.600 ;
        RECT 155.000 66.400 155.800 67.200 ;
        RECT 156.400 66.800 157.200 67.000 ;
        RECT 156.400 66.200 158.800 66.800 ;
        RECT 152.800 64.400 154.400 65.800 ;
        RECT 152.800 63.600 155.600 64.400 ;
        RECT 152.800 62.200 154.400 63.600 ;
        RECT 158.000 62.200 158.800 66.200 ;
        RECT 161.400 64.400 162.000 67.600 ;
        RECT 166.200 67.400 166.800 70.400 ;
        RECT 170.800 71.200 171.400 71.800 ;
        RECT 175.600 71.200 176.200 71.800 ;
        RECT 170.800 70.400 172.000 71.200 ;
        RECT 175.600 70.400 176.800 71.200 ;
        RECT 170.800 67.400 171.400 70.400 ;
        RECT 175.600 67.400 176.200 70.400 ;
        RECT 166.200 66.800 168.400 67.400 ;
        RECT 161.200 62.200 162.000 64.400 ;
        RECT 167.600 62.200 168.400 66.800 ;
        RECT 169.200 66.800 171.400 67.400 ;
        RECT 174.000 66.800 176.200 67.400 ;
        RECT 169.200 62.200 170.000 66.800 ;
        RECT 174.000 62.200 174.800 66.800 ;
        RECT 4.400 55.200 5.200 59.800 ;
        RECT 9.200 55.200 10.000 59.800 ;
        RECT 11.400 58.400 12.200 59.800 ;
        RECT 11.400 57.600 13.200 58.400 ;
        RECT 11.400 56.400 12.200 57.600 ;
        RECT 11.400 55.800 13.200 56.400 ;
        RECT 15.600 55.800 16.400 59.800 ;
        RECT 19.800 58.400 20.600 59.800 ;
        RECT 19.800 57.600 21.200 58.400 ;
        RECT 19.800 56.800 20.600 57.600 ;
        RECT 19.800 55.800 21.200 56.800 ;
        RECT 3.000 54.600 5.200 55.200 ;
        RECT 7.800 54.600 10.000 55.200 ;
        RECT 3.000 51.600 3.600 54.600 ;
        RECT 7.800 51.600 8.400 54.600 ;
        RECT 2.400 50.800 3.600 51.600 ;
        RECT 7.200 50.800 8.400 51.600 ;
        RECT 3.000 50.200 3.600 50.800 ;
        RECT 7.800 50.200 8.400 50.800 ;
        RECT 3.000 49.600 5.200 50.200 ;
        RECT 7.800 49.600 10.000 50.200 ;
        RECT 4.400 42.200 5.200 49.600 ;
        RECT 9.200 42.200 10.000 49.600 ;
        RECT 10.800 48.800 11.600 50.400 ;
        RECT 12.400 42.200 13.200 55.800 ;
        RECT 15.800 55.600 16.400 55.800 ;
        RECT 15.800 55.200 17.600 55.600 ;
        RECT 14.000 54.300 14.800 55.200 ;
        RECT 15.800 55.000 20.000 55.200 ;
        RECT 17.000 54.600 20.000 55.000 ;
        RECT 19.200 54.400 20.000 54.600 ;
        RECT 15.600 54.300 16.400 54.400 ;
        RECT 14.000 53.700 16.400 54.300 ;
        RECT 17.600 53.800 18.400 54.000 ;
        RECT 14.000 53.600 14.800 53.700 ;
        RECT 15.600 52.800 16.400 53.700 ;
        RECT 17.400 53.200 18.400 53.800 ;
        RECT 17.400 52.400 18.000 53.200 ;
        RECT 17.200 51.600 18.000 52.400 ;
        RECT 19.200 51.000 19.800 54.400 ;
        RECT 20.600 52.400 21.200 55.800 ;
        RECT 22.000 55.800 22.800 59.800 ;
        RECT 26.400 56.200 28.000 59.800 ;
        RECT 22.000 55.200 24.400 55.800 ;
        RECT 23.600 55.000 24.400 55.200 ;
        RECT 25.000 54.800 25.800 55.600 ;
        RECT 25.000 54.400 25.600 54.800 ;
        RECT 24.800 53.600 25.600 54.400 ;
        RECT 26.400 52.800 27.000 56.200 ;
        RECT 31.600 55.800 32.400 59.800 ;
        RECT 34.800 57.800 35.600 59.800 ;
        RECT 27.600 55.400 29.200 55.600 ;
        RECT 27.600 54.800 29.600 55.400 ;
        RECT 30.200 55.200 32.400 55.800 ;
        RECT 33.200 56.300 34.000 56.400 ;
        RECT 34.800 56.300 35.400 57.800 ;
        RECT 38.200 56.400 39.000 57.200 ;
        RECT 33.200 55.700 35.500 56.300 ;
        RECT 33.200 55.600 34.000 55.700 ;
        RECT 30.200 55.000 31.000 55.200 ;
        RECT 29.000 54.400 29.600 54.800 ;
        RECT 34.800 54.400 35.400 55.700 ;
        RECT 38.000 55.600 38.800 56.400 ;
        RECT 39.600 55.800 40.400 59.800 ;
        RECT 27.600 53.400 28.400 54.200 ;
        RECT 29.000 53.800 32.400 54.400 ;
        RECT 30.800 53.600 32.400 53.800 ;
        RECT 34.800 53.600 35.600 54.400 ;
        RECT 26.000 52.400 27.000 52.800 ;
        RECT 20.400 51.600 21.200 52.400 ;
        RECT 25.200 52.200 27.000 52.400 ;
        RECT 27.800 52.800 28.400 53.400 ;
        RECT 27.800 52.200 30.400 52.800 ;
        RECT 25.200 51.600 26.600 52.200 ;
        RECT 29.600 52.000 30.400 52.200 ;
        RECT 17.400 50.400 19.800 51.000 ;
        RECT 17.400 46.200 18.000 50.400 ;
        RECT 20.600 50.200 21.200 51.600 ;
        RECT 26.000 50.200 26.600 51.600 ;
        RECT 27.400 51.400 28.200 51.600 ;
        RECT 27.400 50.800 30.800 51.400 ;
        RECT 30.200 50.200 30.800 50.800 ;
        RECT 34.800 50.200 35.400 53.600 ;
        RECT 39.800 52.400 40.400 55.800 ;
        RECT 41.200 52.800 42.000 54.400 ;
        RECT 38.000 52.200 38.800 52.400 ;
        RECT 39.600 52.200 40.400 52.400 ;
        RECT 42.800 52.200 43.600 52.400 ;
        RECT 38.000 51.600 40.400 52.200 ;
        RECT 42.000 51.600 43.600 52.200 ;
        RECT 38.200 50.200 38.800 51.600 ;
        RECT 42.000 51.200 42.800 51.600 ;
        RECT 46.000 50.300 46.800 59.800 ;
        RECT 56.000 54.200 56.800 59.800 ;
        RECT 58.800 56.000 59.600 59.800 ;
        RECT 62.000 56.000 62.800 59.800 ;
        RECT 58.800 55.800 62.800 56.000 ;
        RECT 63.600 55.800 64.400 59.800 ;
        RECT 67.800 58.400 68.600 59.800 ;
        RECT 67.800 57.600 69.200 58.400 ;
        RECT 67.800 56.400 68.600 57.600 ;
        RECT 66.800 55.800 68.600 56.400 ;
        RECT 59.000 55.400 62.600 55.800 ;
        RECT 63.600 54.400 64.200 55.800 ;
        RECT 56.000 53.800 57.800 54.200 ;
        RECT 56.200 53.600 57.800 53.800 ;
        RECT 54.000 51.600 55.600 52.400 ;
        RECT 57.200 52.300 57.800 53.600 ;
        RECT 61.800 53.600 64.400 54.400 ;
        RECT 60.400 52.300 61.200 53.200 ;
        RECT 57.200 51.700 61.200 52.300 ;
        RECT 52.400 50.300 53.200 51.200 ;
        RECT 17.200 42.200 18.000 46.200 ;
        RECT 20.400 42.200 21.200 50.200 ;
        RECT 22.000 49.600 24.400 50.200 ;
        RECT 26.000 49.600 28.000 50.200 ;
        RECT 22.000 42.200 22.800 49.600 ;
        RECT 23.600 49.400 24.400 49.600 ;
        RECT 26.400 44.400 28.000 49.600 ;
        RECT 30.200 49.600 32.400 50.200 ;
        RECT 30.200 49.400 31.000 49.600 ;
        RECT 25.200 43.600 28.000 44.400 ;
        RECT 26.400 42.200 28.000 43.600 ;
        RECT 31.600 42.200 32.400 49.600 ;
        RECT 33.800 49.400 35.600 50.200 ;
        RECT 33.800 42.200 34.600 49.400 ;
        RECT 38.000 42.200 38.800 50.200 ;
        RECT 39.600 49.600 43.600 50.200 ;
        RECT 39.600 42.200 40.400 49.600 ;
        RECT 42.800 42.200 43.600 49.600 ;
        RECT 46.000 49.700 53.200 50.300 ;
        RECT 46.000 42.200 46.800 49.700 ;
        RECT 52.400 49.600 53.200 49.700 ;
        RECT 57.200 50.400 57.800 51.700 ;
        RECT 60.400 51.600 61.200 51.700 ;
        RECT 61.800 52.300 62.400 53.600 ;
        RECT 65.200 52.300 66.000 52.400 ;
        RECT 61.800 51.700 66.000 52.300 ;
        RECT 57.200 49.600 58.000 50.400 ;
        RECT 61.800 50.200 62.400 51.700 ;
        RECT 65.200 51.600 66.000 51.700 ;
        RECT 63.600 50.200 64.400 50.400 ;
        RECT 61.400 49.600 62.400 50.200 ;
        RECT 63.000 49.600 64.400 50.200 ;
        RECT 55.600 47.600 56.400 49.200 ;
        RECT 57.200 47.000 57.800 49.600 ;
        RECT 54.200 46.400 57.800 47.000 ;
        RECT 54.000 42.200 54.800 46.400 ;
        RECT 57.200 46.200 57.800 46.400 ;
        RECT 57.200 42.200 58.000 46.200 ;
        RECT 61.400 42.200 62.200 49.600 ;
        RECT 63.000 48.400 63.600 49.600 ;
        RECT 62.800 47.600 63.600 48.400 ;
        RECT 66.800 42.200 67.600 55.800 ;
        RECT 68.400 48.800 69.200 50.400 ;
        RECT 70.000 42.200 70.800 59.800 ;
        RECT 74.800 57.800 75.600 59.800 ;
        RECT 71.600 56.300 72.400 57.200 ;
        RECT 73.200 56.300 74.000 56.400 ;
        RECT 71.600 55.700 74.000 56.300 ;
        RECT 71.600 55.600 72.400 55.700 ;
        RECT 73.200 55.600 74.000 55.700 ;
        RECT 74.800 54.400 75.400 57.800 ;
        RECT 76.400 55.600 77.200 57.200 ;
        RECT 74.800 53.600 75.600 54.400 ;
        RECT 74.800 52.400 75.400 53.600 ;
        RECT 78.000 52.400 78.800 59.800 ;
        RECT 81.200 55.200 82.000 59.800 ;
        RECT 83.400 58.400 84.200 59.800 ;
        RECT 83.400 57.600 85.200 58.400 ;
        RECT 92.400 57.800 93.200 59.800 ;
        RECT 95.600 58.400 96.400 59.800 ;
        RECT 92.000 57.600 93.200 57.800 ;
        RECT 95.400 57.600 96.400 58.400 ;
        RECT 83.400 56.400 84.200 57.600 ;
        RECT 92.000 57.000 96.000 57.600 ;
        RECT 83.400 55.800 85.200 56.400 ;
        RECT 79.800 54.600 82.000 55.200 ;
        RECT 73.200 50.800 74.000 52.400 ;
        RECT 74.800 51.600 75.600 52.400 ;
        RECT 74.800 50.200 75.400 51.600 ;
        RECT 78.000 50.200 78.600 52.400 ;
        RECT 79.800 51.600 80.400 54.600 ;
        RECT 81.200 51.600 82.000 53.200 ;
        RECT 79.200 50.800 80.400 51.600 ;
        RECT 79.800 50.200 80.400 50.800 ;
        RECT 73.800 49.400 75.600 50.200 ;
        RECT 73.800 42.200 74.600 49.400 ;
        RECT 78.000 42.200 78.800 50.200 ;
        RECT 79.800 49.600 82.000 50.200 ;
        RECT 81.200 42.200 82.000 49.600 ;
        RECT 82.800 48.800 83.600 50.400 ;
        RECT 84.400 42.200 85.200 55.800 ;
        RECT 86.000 53.600 86.800 55.200 ;
        RECT 92.000 50.400 92.600 57.000 ;
        RECT 101.000 56.400 101.800 59.800 ;
        RECT 105.800 56.800 106.600 59.800 ;
        RECT 96.200 55.600 98.000 56.400 ;
        RECT 101.000 55.800 102.800 56.400 ;
        RECT 94.800 54.300 96.400 54.400 ;
        RECT 98.800 54.300 99.600 54.400 ;
        RECT 94.800 53.700 99.600 54.300 ;
        RECT 94.800 53.600 96.400 53.700 ;
        RECT 98.800 53.600 99.600 53.700 ;
        RECT 93.200 52.300 94.800 52.400 ;
        RECT 97.200 52.300 98.000 52.400 ;
        RECT 93.200 51.700 98.000 52.300 ;
        RECT 93.200 51.600 94.800 51.700 ;
        RECT 97.200 51.600 98.000 51.700 ;
        RECT 89.200 49.800 92.600 50.400 ;
        RECT 89.200 49.600 90.000 49.800 ;
        RECT 89.400 49.000 90.000 49.600 ;
        RECT 91.000 49.000 94.600 49.200 ;
        RECT 87.600 43.000 88.400 49.000 ;
        RECT 89.200 43.400 90.000 49.000 ;
        RECT 90.800 48.600 94.600 49.000 ;
        RECT 87.800 42.800 88.400 43.000 ;
        RECT 90.800 43.000 91.600 48.600 ;
        RECT 94.000 48.200 94.600 48.600 ;
        RECT 95.800 48.800 99.400 49.400 ;
        RECT 100.400 48.800 101.200 50.400 ;
        RECT 95.800 48.200 96.400 48.800 ;
        RECT 90.800 42.800 91.400 43.000 ;
        RECT 87.800 42.200 91.400 42.800 ;
        RECT 92.400 42.800 93.200 48.000 ;
        RECT 94.000 43.400 94.800 48.200 ;
        RECT 95.600 42.800 96.400 48.200 ;
        RECT 92.400 42.200 96.400 42.800 ;
        RECT 98.800 48.200 99.400 48.800 ;
        RECT 98.800 42.200 99.600 48.200 ;
        RECT 102.000 42.200 102.800 55.800 ;
        RECT 105.200 55.800 106.600 56.800 ;
        RECT 110.000 55.800 110.800 59.800 ;
        RECT 112.200 58.400 113.000 59.800 ;
        RECT 111.600 57.600 113.000 58.400 ;
        RECT 112.200 56.400 113.000 57.600 ;
        RECT 117.000 56.400 117.800 59.800 ;
        RECT 112.200 55.800 114.000 56.400 ;
        RECT 117.000 55.800 118.800 56.400 ;
        RECT 103.600 53.600 104.400 55.200 ;
        RECT 103.700 52.400 104.300 53.600 ;
        RECT 105.200 52.400 105.800 55.800 ;
        RECT 110.000 55.600 110.600 55.800 ;
        RECT 108.800 55.200 110.600 55.600 ;
        RECT 106.400 55.000 110.600 55.200 ;
        RECT 106.400 54.600 109.400 55.000 ;
        RECT 106.400 54.400 107.200 54.600 ;
        RECT 103.600 52.300 104.400 52.400 ;
        RECT 105.200 52.300 106.000 52.400 ;
        RECT 103.600 51.700 106.000 52.300 ;
        RECT 103.600 51.600 104.400 51.700 ;
        RECT 105.200 51.600 106.000 51.700 ;
        RECT 105.200 50.200 105.800 51.600 ;
        RECT 106.600 51.000 107.200 54.400 ;
        RECT 108.000 53.800 108.800 54.000 ;
        RECT 108.000 53.200 109.000 53.800 ;
        RECT 108.400 52.400 109.000 53.200 ;
        RECT 110.000 52.800 110.800 54.400 ;
        RECT 108.400 51.600 109.200 52.400 ;
        RECT 106.600 50.400 109.000 51.000 ;
        RECT 105.200 42.200 106.000 50.200 ;
        RECT 108.400 46.200 109.000 50.400 ;
        RECT 111.600 48.800 112.400 50.400 ;
        RECT 108.400 42.200 109.200 46.200 ;
        RECT 113.200 42.200 114.000 55.800 ;
        RECT 114.800 53.600 115.600 55.200 ;
        RECT 116.400 48.800 117.200 50.400 ;
        RECT 118.000 42.200 118.800 55.800 ;
        RECT 119.600 53.600 120.400 55.200 ;
        RECT 121.200 52.400 122.000 59.800 ;
        RECT 124.400 55.200 125.200 59.800 ;
        RECT 123.000 54.600 125.200 55.200 ;
        RECT 130.800 55.200 131.600 59.800 ;
        RECT 130.800 54.600 133.000 55.200 ;
        RECT 121.200 50.200 121.800 52.400 ;
        RECT 123.000 51.600 123.600 54.600 ;
        RECT 124.400 52.300 125.200 53.200 ;
        RECT 130.800 52.300 131.600 53.200 ;
        RECT 124.400 51.700 131.600 52.300 ;
        RECT 124.400 51.600 125.200 51.700 ;
        RECT 130.800 51.600 131.600 51.700 ;
        RECT 132.400 51.600 133.000 54.600 ;
        RECT 134.000 52.400 134.800 59.800 ;
        RECT 137.200 57.800 138.000 59.800 ;
        RECT 137.200 54.400 137.800 57.800 ;
        RECT 138.800 55.600 139.600 57.200 ;
        RECT 140.400 55.800 141.200 59.800 ;
        RECT 144.800 56.200 146.400 59.800 ;
        RECT 140.400 55.200 143.000 55.800 ;
        RECT 142.200 55.000 143.000 55.200 ;
        RECT 143.600 54.800 145.200 55.600 ;
        RECT 137.200 54.300 138.000 54.400 ;
        RECT 138.800 54.300 139.600 54.400 ;
        RECT 137.200 53.700 139.600 54.300 ;
        RECT 137.200 53.600 138.000 53.700 ;
        RECT 138.800 53.600 139.600 53.700 ;
        RECT 140.400 54.200 142.000 54.400 ;
        RECT 145.800 54.200 146.400 56.200 ;
        RECT 150.000 55.800 150.800 59.800 ;
        RECT 154.800 58.400 155.600 59.800 ;
        RECT 154.800 57.800 155.800 58.400 ;
        RECT 155.200 57.600 155.800 57.800 ;
        RECT 158.000 57.800 158.800 59.800 ;
        RECT 158.000 57.600 159.200 57.800 ;
        RECT 155.200 57.000 159.200 57.600 ;
        RECT 147.000 54.800 147.800 55.600 ;
        RECT 148.400 55.200 150.800 55.800 ;
        RECT 153.200 56.300 155.000 56.400 ;
        RECT 156.400 56.300 157.200 56.400 ;
        RECT 153.200 55.700 157.200 56.300 ;
        RECT 153.200 55.600 155.000 55.700 ;
        RECT 156.400 55.600 157.200 55.700 ;
        RECT 148.400 55.000 149.200 55.200 ;
        RECT 140.400 54.000 142.600 54.200 ;
        RECT 140.400 53.600 144.800 54.000 ;
        RECT 122.400 50.800 123.600 51.600 ;
        RECT 123.000 50.200 123.600 50.800 ;
        RECT 132.400 50.800 133.600 51.600 ;
        RECT 132.400 50.200 133.000 50.800 ;
        RECT 134.200 50.200 134.800 52.400 ;
        RECT 135.600 50.800 136.400 52.400 ;
        RECT 137.200 50.200 137.800 53.600 ;
        RECT 142.000 53.400 144.800 53.600 ;
        RECT 144.000 53.200 144.800 53.400 ;
        RECT 145.400 53.600 146.400 54.200 ;
        RECT 147.200 54.400 147.800 54.800 ;
        RECT 147.200 53.600 148.000 54.400 ;
        RECT 154.800 53.600 156.400 54.400 ;
        RECT 145.400 52.400 146.000 53.600 ;
        RECT 142.600 52.200 143.400 52.400 ;
        RECT 142.600 51.600 144.200 52.200 ;
        RECT 145.200 51.600 146.000 52.400 ;
        RECT 156.400 51.600 158.000 52.400 ;
        RECT 143.400 51.400 144.200 51.600 ;
        RECT 145.400 50.200 146.000 51.600 ;
        RECT 158.600 50.400 159.200 57.000 ;
        RECT 164.400 55.200 165.200 59.800 ;
        RECT 169.200 55.200 170.000 59.800 ;
        RECT 175.600 57.600 176.400 59.800 ;
        RECT 164.400 54.600 166.600 55.200 ;
        RECT 169.200 54.600 171.400 55.200 ;
        RECT 164.400 51.600 165.200 53.200 ;
        RECT 166.000 51.600 166.600 54.600 ;
        RECT 169.200 51.600 170.000 53.200 ;
        RECT 170.800 51.600 171.400 54.600 ;
        RECT 175.800 54.400 176.400 57.600 ;
        RECT 175.600 53.600 176.400 54.400 ;
        RECT 166.000 50.800 167.200 51.600 ;
        RECT 170.800 50.800 172.000 51.600 ;
        RECT 121.200 42.200 122.000 50.200 ;
        RECT 123.000 49.600 125.200 50.200 ;
        RECT 124.400 42.200 125.200 49.600 ;
        RECT 130.800 49.600 133.000 50.200 ;
        RECT 130.800 42.200 131.600 49.600 ;
        RECT 134.000 42.200 134.800 50.200 ;
        RECT 136.200 49.400 138.000 50.200 ;
        RECT 140.400 49.600 143.000 50.200 ;
        RECT 136.200 42.200 137.000 49.400 ;
        RECT 140.400 42.200 141.200 49.600 ;
        RECT 142.200 49.400 143.000 49.600 ;
        RECT 144.800 44.400 146.400 50.200 ;
        RECT 148.400 49.600 150.800 50.200 ;
        RECT 158.600 49.800 162.000 50.400 ;
        RECT 166.000 50.200 166.600 50.800 ;
        RECT 170.800 50.200 171.400 50.800 ;
        RECT 175.800 50.200 176.400 53.600 ;
        RECT 148.400 49.400 149.200 49.600 ;
        RECT 143.600 43.600 146.400 44.400 ;
        RECT 144.800 42.200 146.400 43.600 ;
        RECT 150.000 42.200 150.800 49.600 ;
        RECT 161.200 49.600 162.000 49.800 ;
        RECT 164.400 49.600 166.600 50.200 ;
        RECT 169.200 49.600 171.400 50.200 ;
        RECT 151.800 48.800 155.400 49.400 ;
        RECT 151.800 48.200 152.400 48.800 ;
        RECT 151.600 42.200 152.400 48.200 ;
        RECT 154.800 48.200 155.400 48.800 ;
        RECT 156.600 49.000 160.200 49.200 ;
        RECT 161.200 49.000 161.800 49.600 ;
        RECT 156.600 48.600 160.400 49.000 ;
        RECT 156.600 48.200 157.200 48.600 ;
        RECT 154.800 42.800 155.600 48.200 ;
        RECT 156.400 43.400 157.200 48.200 ;
        RECT 158.000 42.800 158.800 48.000 ;
        RECT 159.600 43.000 160.400 48.600 ;
        RECT 161.200 43.400 162.000 49.000 ;
        RECT 154.800 42.200 158.800 42.800 ;
        RECT 159.800 42.800 160.400 43.000 ;
        RECT 162.800 43.000 163.600 49.000 ;
        RECT 162.800 42.800 163.400 43.000 ;
        RECT 159.800 42.200 163.400 42.800 ;
        RECT 164.400 42.200 165.200 49.600 ;
        RECT 169.200 42.200 170.000 49.600 ;
        RECT 175.600 49.400 177.400 50.200 ;
        RECT 176.600 44.400 177.400 49.400 ;
        RECT 175.600 43.600 177.400 44.400 ;
        RECT 176.600 42.200 177.400 43.600 ;
        RECT 1.400 39.200 5.000 39.800 ;
        RECT 1.400 39.000 2.000 39.200 ;
        RECT 1.200 33.000 2.000 39.000 ;
        RECT 4.400 39.000 5.000 39.200 ;
        RECT 6.000 39.200 10.000 39.800 ;
        RECT 2.800 33.000 3.600 38.600 ;
        RECT 4.400 33.400 5.200 39.000 ;
        RECT 6.000 34.000 6.800 39.200 ;
        RECT 7.600 33.800 8.400 38.600 ;
        RECT 9.200 33.800 10.000 39.200 ;
        RECT 7.600 33.400 8.200 33.800 ;
        RECT 4.400 33.000 8.200 33.400 ;
        RECT 3.000 32.400 3.600 33.000 ;
        RECT 4.600 32.800 8.200 33.000 ;
        RECT 9.400 33.200 10.000 33.800 ;
        RECT 12.400 33.800 13.200 39.800 ;
        RECT 12.400 33.200 13.000 33.800 ;
        RECT 9.400 32.600 13.000 33.200 ;
        RECT 14.600 32.400 15.400 39.800 ;
        RECT 2.800 32.200 3.600 32.400 ;
        RECT 2.800 31.600 6.200 32.200 ;
        RECT 5.600 25.000 6.200 31.600 ;
        RECT 14.000 31.800 15.400 32.400 ;
        RECT 14.000 30.400 14.600 31.800 ;
        RECT 18.800 31.200 19.600 39.800 ;
        RECT 23.000 38.400 23.800 39.800 ;
        RECT 22.000 37.600 23.800 38.400 ;
        RECT 23.000 32.400 23.800 37.600 ;
        RECT 24.400 33.600 25.200 34.400 ;
        RECT 24.600 32.400 25.200 33.600 ;
        RECT 23.000 31.800 24.000 32.400 ;
        RECT 24.600 31.800 26.000 32.400 ;
        RECT 15.600 30.800 19.600 31.200 ;
        RECT 15.400 30.600 19.600 30.800 ;
        RECT 6.800 29.600 8.400 30.400 ;
        RECT 14.000 29.600 14.800 30.400 ;
        RECT 15.400 30.000 16.200 30.600 ;
        RECT 8.400 27.600 10.000 28.400 ;
        RECT 9.800 25.600 11.600 26.400 ;
        RECT 14.000 26.200 14.600 29.600 ;
        RECT 15.400 27.000 16.000 30.000 ;
        RECT 16.800 28.400 17.600 29.200 ;
        RECT 22.000 28.800 22.800 30.400 ;
        RECT 23.400 28.400 24.000 31.800 ;
        RECT 25.200 31.600 26.000 31.800 ;
        RECT 17.000 27.600 18.000 28.400 ;
        RECT 20.400 28.300 21.200 28.400 ;
        RECT 18.900 28.200 21.200 28.300 ;
        RECT 18.900 27.700 22.000 28.200 ;
        RECT 15.400 26.400 17.800 27.000 ;
        RECT 18.900 26.400 19.500 27.700 ;
        RECT 20.400 27.600 22.000 27.700 ;
        RECT 23.400 27.600 26.000 28.400 ;
        RECT 21.200 27.200 22.000 27.600 ;
        RECT 5.600 24.400 9.600 25.000 ;
        RECT 4.400 23.600 6.800 24.400 ;
        RECT 9.000 24.200 9.600 24.400 ;
        RECT 9.000 23.600 10.000 24.200 ;
        RECT 6.000 22.200 6.800 23.600 ;
        RECT 9.200 22.200 10.000 23.600 ;
        RECT 14.000 22.200 14.800 26.200 ;
        RECT 17.200 24.200 17.800 26.400 ;
        RECT 18.800 24.800 19.600 26.400 ;
        RECT 20.600 26.200 24.200 26.600 ;
        RECT 25.200 26.200 25.800 27.600 ;
        RECT 20.400 26.000 24.400 26.200 ;
        RECT 17.200 22.200 18.000 24.200 ;
        RECT 20.400 22.200 21.200 26.000 ;
        RECT 23.600 22.200 24.400 26.000 ;
        RECT 25.200 22.200 26.000 26.200 ;
        RECT 26.800 22.200 27.600 39.800 ;
        RECT 30.000 35.800 30.800 39.800 ;
        RECT 30.200 35.600 30.800 35.800 ;
        RECT 33.200 35.800 34.000 39.800 ;
        RECT 33.200 35.600 33.800 35.800 ;
        RECT 30.200 35.000 33.800 35.600 ;
        RECT 30.200 32.400 30.800 35.000 ;
        RECT 31.600 32.800 32.400 34.400 ;
        RECT 30.000 31.600 30.800 32.400 ;
        RECT 30.200 28.400 30.800 31.600 ;
        RECT 34.800 30.800 35.600 32.400 ;
        RECT 36.400 31.800 37.200 39.800 ;
        RECT 38.000 32.400 38.800 39.800 ;
        RECT 41.200 32.400 42.000 39.800 ;
        RECT 38.000 31.800 42.000 32.400 ;
        RECT 42.800 32.400 43.600 39.800 ;
        RECT 44.200 32.400 45.000 32.600 ;
        RECT 42.800 31.800 45.000 32.400 ;
        RECT 47.200 32.400 48.800 39.800 ;
        RECT 50.800 32.400 51.600 32.600 ;
        RECT 52.400 32.400 53.200 39.800 ;
        RECT 59.000 39.200 62.600 39.800 ;
        RECT 59.000 39.000 59.600 39.200 ;
        RECT 58.800 33.000 59.600 39.000 ;
        RECT 62.000 39.000 62.600 39.200 ;
        RECT 63.600 39.200 67.600 39.800 ;
        RECT 60.400 33.000 61.200 38.600 ;
        RECT 62.000 33.400 62.800 39.000 ;
        RECT 63.600 34.000 64.400 39.200 ;
        RECT 65.200 33.800 66.000 38.600 ;
        RECT 66.800 33.800 67.600 39.200 ;
        RECT 65.200 33.400 65.800 33.800 ;
        RECT 62.000 33.000 65.800 33.400 ;
        RECT 60.600 32.400 61.200 33.000 ;
        RECT 62.200 32.800 65.800 33.000 ;
        RECT 67.000 33.200 67.600 33.800 ;
        RECT 70.000 33.800 70.800 39.800 ;
        RECT 70.000 33.200 70.600 33.800 ;
        RECT 67.000 32.600 70.600 33.200 ;
        RECT 47.200 31.800 49.200 32.400 ;
        RECT 50.800 31.800 53.200 32.400 ;
        RECT 60.400 32.200 61.200 32.400 ;
        RECT 36.600 30.400 37.200 31.800 ;
        RECT 44.400 31.200 45.000 31.800 ;
        RECT 40.400 30.400 41.200 30.800 ;
        RECT 44.400 30.600 47.800 31.200 ;
        RECT 47.000 30.400 47.800 30.600 ;
        RECT 48.600 30.400 49.200 31.800 ;
        RECT 60.400 31.600 63.800 32.200 ;
        RECT 36.400 29.800 38.800 30.400 ;
        RECT 40.400 29.800 42.000 30.400 ;
        RECT 36.400 29.600 37.200 29.800 ;
        RECT 38.200 28.400 38.800 29.800 ;
        RECT 41.200 29.600 42.000 29.800 ;
        RECT 44.800 29.800 45.600 30.000 ;
        RECT 48.600 29.800 50.000 30.400 ;
        RECT 44.800 29.200 47.400 29.800 ;
        RECT 30.200 28.200 31.800 28.400 ;
        RECT 30.200 27.800 32.000 28.200 ;
        RECT 28.400 26.300 29.200 26.400 ;
        RECT 31.200 26.300 32.000 27.800 ;
        RECT 38.000 27.600 38.800 28.400 ;
        RECT 39.600 27.600 40.400 29.200 ;
        RECT 46.800 28.600 47.400 29.200 ;
        RECT 48.200 29.600 50.000 29.800 ;
        RECT 48.200 29.200 49.200 29.600 ;
        RECT 42.800 28.200 44.400 28.400 ;
        RECT 42.800 27.600 46.200 28.200 ;
        RECT 46.800 27.800 47.600 28.600 ;
        RECT 28.400 25.700 32.000 26.300 ;
        RECT 38.200 26.200 38.800 27.600 ;
        RECT 45.600 27.200 46.200 27.600 ;
        RECT 44.200 26.800 45.000 27.000 ;
        RECT 28.400 24.800 29.200 25.700 ;
        RECT 31.200 22.200 32.000 25.700 ;
        RECT 38.000 22.200 38.800 26.200 ;
        RECT 42.800 26.200 45.000 26.800 ;
        RECT 45.600 26.600 47.600 27.200 ;
        RECT 46.000 26.400 47.600 26.600 ;
        RECT 42.800 22.200 43.600 26.200 ;
        RECT 48.200 25.800 48.800 29.200 ;
        RECT 49.600 27.600 50.400 28.400 ;
        RECT 49.600 27.200 50.200 27.600 ;
        RECT 49.400 26.400 50.200 27.200 ;
        RECT 50.800 26.800 51.600 27.000 ;
        RECT 50.800 26.200 53.200 26.800 ;
        RECT 47.200 24.400 48.800 25.800 ;
        RECT 46.000 23.600 48.800 24.400 ;
        RECT 47.200 22.200 48.800 23.600 ;
        RECT 52.400 22.200 53.200 26.200 ;
        RECT 63.200 25.000 63.800 31.600 ;
        RECT 64.400 29.600 66.000 30.400 ;
        RECT 73.200 30.300 74.000 39.800 ;
        RECT 77.400 32.400 78.200 39.800 ;
        RECT 78.800 33.600 79.600 34.400 ;
        RECT 79.000 32.400 79.600 33.600 ;
        RECT 81.200 32.400 82.000 39.800 ;
        RECT 82.800 32.400 83.600 32.600 ;
        RECT 85.600 32.400 87.200 39.800 ;
        RECT 76.400 31.600 78.400 32.400 ;
        RECT 79.000 31.800 80.400 32.400 ;
        RECT 81.200 31.800 83.600 32.400 ;
        RECT 85.200 31.800 87.200 32.400 ;
        RECT 89.400 32.400 90.200 32.600 ;
        RECT 90.800 32.400 91.600 39.800 ;
        RECT 95.600 32.400 96.400 39.800 ;
        RECT 89.400 31.800 91.600 32.400 ;
        RECT 94.200 31.800 96.400 32.400 ;
        RECT 79.600 31.600 80.400 31.800 ;
        RECT 76.400 30.300 77.200 30.400 ;
        RECT 73.200 29.700 77.200 30.300 ;
        RECT 66.000 28.300 67.600 28.400 ;
        RECT 70.000 28.300 70.800 28.400 ;
        RECT 66.000 27.700 70.800 28.300 ;
        RECT 66.000 27.600 67.600 27.700 ;
        RECT 70.000 27.600 70.800 27.700 ;
        RECT 67.400 25.600 69.200 26.400 ;
        RECT 63.200 24.400 67.200 25.000 ;
        RECT 57.200 24.300 58.000 24.400 ;
        RECT 63.200 24.300 64.400 24.400 ;
        RECT 57.200 23.700 64.400 24.300 ;
        RECT 57.200 23.600 58.000 23.700 ;
        RECT 63.600 22.200 64.400 23.700 ;
        RECT 66.600 24.200 67.200 24.400 ;
        RECT 66.600 23.600 67.600 24.200 ;
        RECT 66.800 22.200 67.600 23.600 ;
        RECT 73.200 22.200 74.000 29.700 ;
        RECT 76.400 28.800 77.200 29.700 ;
        RECT 77.800 28.400 78.400 31.600 ;
        RECT 85.200 30.400 85.800 31.800 ;
        RECT 89.400 31.200 90.000 31.800 ;
        RECT 94.200 31.200 94.800 31.800 ;
        RECT 86.600 30.600 90.000 31.200 ;
        RECT 86.600 30.400 87.400 30.600 ;
        RECT 93.600 30.400 94.800 31.200 ;
        RECT 84.400 29.800 85.800 30.400 ;
        RECT 88.800 29.800 89.600 30.000 ;
        RECT 84.400 29.600 86.200 29.800 ;
        RECT 85.200 29.200 86.200 29.600 ;
        RECT 74.800 28.200 75.600 28.400 ;
        RECT 74.800 27.600 76.400 28.200 ;
        RECT 77.800 27.600 80.400 28.400 ;
        RECT 81.200 27.600 82.800 28.400 ;
        RECT 84.000 27.600 84.800 28.400 ;
        RECT 75.600 27.200 76.400 27.600 ;
        RECT 75.000 26.200 78.600 26.600 ;
        RECT 79.600 26.200 80.200 27.600 ;
        RECT 84.200 27.200 84.800 27.600 ;
        RECT 82.800 26.800 83.600 27.000 ;
        RECT 81.200 26.200 83.600 26.800 ;
        RECT 84.200 26.400 85.000 27.200 ;
        RECT 74.800 26.000 78.800 26.200 ;
        RECT 74.800 22.200 75.600 26.000 ;
        RECT 78.000 22.200 78.800 26.000 ;
        RECT 79.600 22.200 80.400 26.200 ;
        RECT 81.200 22.200 82.000 26.200 ;
        RECT 85.600 25.800 86.200 29.200 ;
        RECT 87.000 29.200 89.600 29.800 ;
        RECT 87.000 28.600 87.600 29.200 ;
        RECT 86.800 27.800 87.600 28.600 ;
        RECT 90.000 28.200 91.600 28.400 ;
        RECT 88.200 27.600 91.600 28.200 ;
        RECT 88.200 27.200 88.800 27.600 ;
        RECT 86.800 26.600 88.800 27.200 ;
        RECT 94.200 27.400 94.800 30.400 ;
        RECT 95.600 28.800 96.400 30.400 ;
        RECT 98.800 28.300 99.600 39.800 ;
        RECT 103.000 32.400 103.800 39.800 ;
        RECT 104.400 33.600 105.200 34.400 ;
        RECT 104.600 32.400 105.200 33.600 ;
        RECT 109.400 32.400 110.200 39.800 ;
        RECT 110.800 33.600 111.600 34.400 ;
        RECT 111.000 32.400 111.600 33.600 ;
        RECT 103.000 31.800 104.000 32.400 ;
        RECT 104.600 31.800 106.000 32.400 ;
        RECT 109.400 31.800 110.400 32.400 ;
        RECT 111.000 31.800 112.400 32.400 ;
        RECT 103.400 30.400 104.000 31.800 ;
        RECT 105.200 31.600 106.000 31.800 ;
        RECT 102.000 28.800 102.800 30.400 ;
        RECT 103.400 29.600 104.400 30.400 ;
        RECT 106.800 30.300 107.600 30.400 ;
        RECT 108.400 30.300 109.200 30.400 ;
        RECT 106.800 29.700 109.200 30.300 ;
        RECT 106.800 29.600 107.600 29.700 ;
        RECT 103.400 28.400 104.000 29.600 ;
        RECT 108.400 28.800 109.200 29.700 ;
        RECT 109.800 28.400 110.400 31.800 ;
        RECT 111.600 31.600 112.400 31.800 ;
        RECT 100.400 28.300 101.200 28.400 ;
        RECT 98.800 28.200 101.200 28.300 ;
        RECT 98.800 27.700 102.000 28.200 ;
        RECT 89.400 26.800 90.200 27.000 ;
        RECT 94.200 26.800 96.400 27.400 ;
        RECT 86.800 26.400 88.400 26.600 ;
        RECT 89.400 26.200 91.600 26.800 ;
        RECT 85.600 24.400 87.200 25.800 ;
        RECT 85.600 23.600 88.400 24.400 ;
        RECT 85.600 22.200 87.200 23.600 ;
        RECT 90.800 22.200 91.600 26.200 ;
        RECT 95.600 22.200 96.400 26.800 ;
        RECT 97.200 24.800 98.000 26.400 ;
        RECT 98.800 22.200 99.600 27.700 ;
        RECT 100.400 27.600 102.000 27.700 ;
        RECT 103.400 27.600 106.000 28.400 ;
        RECT 109.800 27.600 112.400 28.400 ;
        RECT 101.200 27.200 102.000 27.600 ;
        RECT 100.600 26.200 104.200 26.600 ;
        RECT 105.200 26.200 105.800 27.600 ;
        RECT 107.000 26.200 110.600 26.600 ;
        RECT 111.600 26.200 112.200 27.600 ;
        RECT 113.200 26.800 114.000 28.400 ;
        RECT 114.800 26.200 115.600 39.800 ;
        RECT 120.600 38.400 121.400 39.800 ;
        RECT 119.600 37.600 121.400 38.400 ;
        RECT 116.400 31.600 117.200 33.200 ;
        RECT 120.600 32.600 121.400 37.600 ;
        RECT 119.600 31.800 121.400 32.600 ;
        RECT 130.200 32.400 131.000 39.800 ;
        RECT 134.200 39.200 137.800 39.800 ;
        RECT 134.200 39.000 134.800 39.200 ;
        RECT 131.600 33.600 132.400 34.400 ;
        RECT 131.800 32.400 132.400 33.600 ;
        RECT 134.000 33.000 134.800 39.000 ;
        RECT 137.200 39.000 137.800 39.200 ;
        RECT 138.800 39.200 142.800 39.800 ;
        RECT 135.600 33.000 136.400 38.600 ;
        RECT 137.200 33.400 138.000 39.000 ;
        RECT 138.800 34.000 139.600 39.200 ;
        RECT 140.400 33.800 141.200 38.600 ;
        RECT 142.000 33.800 142.800 39.200 ;
        RECT 140.400 33.400 141.000 33.800 ;
        RECT 137.200 33.000 141.000 33.400 ;
        RECT 135.800 32.400 136.400 33.000 ;
        RECT 137.400 32.800 141.000 33.000 ;
        RECT 142.200 33.200 142.800 33.800 ;
        RECT 145.200 33.800 146.000 39.800 ;
        RECT 145.200 33.200 145.800 33.800 ;
        RECT 142.200 32.600 145.800 33.200 ;
        RECT 130.200 31.800 131.200 32.400 ;
        RECT 131.800 31.800 133.200 32.400 ;
        RECT 119.800 28.400 120.400 31.800 ;
        RECT 129.200 28.800 130.000 30.400 ;
        RECT 119.600 27.600 120.400 28.400 ;
        RECT 130.600 28.400 131.200 31.800 ;
        RECT 132.400 31.600 133.200 31.800 ;
        RECT 135.600 32.200 136.400 32.400 ;
        RECT 146.800 32.400 147.600 39.800 ;
        RECT 148.600 32.400 149.400 32.600 ;
        RECT 135.600 31.600 139.000 32.200 ;
        RECT 146.800 31.800 149.400 32.400 ;
        RECT 151.200 31.800 152.800 39.800 ;
        RECT 154.800 32.400 155.600 32.600 ;
        RECT 156.400 32.400 157.200 39.800 ;
        RECT 158.000 33.800 158.800 39.800 ;
        RECT 158.200 33.200 158.800 33.800 ;
        RECT 161.200 39.200 165.200 39.800 ;
        RECT 161.200 33.800 162.000 39.200 ;
        RECT 162.800 33.800 163.600 38.600 ;
        RECT 164.400 34.000 165.200 39.200 ;
        RECT 166.200 39.200 169.800 39.800 ;
        RECT 166.200 39.000 166.800 39.200 ;
        RECT 161.200 33.200 161.800 33.800 ;
        RECT 158.200 32.600 161.800 33.200 ;
        RECT 163.000 33.400 163.600 33.800 ;
        RECT 166.000 33.400 166.800 39.000 ;
        RECT 169.200 39.000 169.800 39.200 ;
        RECT 163.000 33.000 166.800 33.400 ;
        RECT 167.600 33.000 168.400 38.600 ;
        RECT 169.200 33.000 170.000 39.000 ;
        RECT 163.000 32.800 166.600 33.000 ;
        RECT 154.800 31.800 157.200 32.400 ;
        RECT 167.600 32.400 168.200 33.000 ;
        RECT 170.800 32.400 171.600 39.800 ;
        RECT 167.600 32.200 168.400 32.400 ;
        RECT 130.600 28.300 133.200 28.400 ;
        RECT 135.600 28.300 136.400 28.400 ;
        RECT 130.600 27.700 136.400 28.300 ;
        RECT 130.600 27.600 133.200 27.700 ;
        RECT 135.600 27.600 136.400 27.700 ;
        RECT 100.400 26.000 104.400 26.200 ;
        RECT 100.400 22.200 101.200 26.000 ;
        RECT 103.600 22.200 104.400 26.000 ;
        RECT 105.200 22.200 106.000 26.200 ;
        RECT 106.800 26.000 110.800 26.200 ;
        RECT 106.800 22.200 107.600 26.000 ;
        RECT 110.000 22.200 110.800 26.000 ;
        RECT 111.600 22.200 112.400 26.200 ;
        RECT 114.800 25.600 116.600 26.200 ;
        RECT 115.800 24.400 116.600 25.600 ;
        RECT 114.800 23.600 116.600 24.400 ;
        RECT 119.800 24.200 120.400 27.600 ;
        RECT 127.800 26.200 131.400 26.600 ;
        RECT 132.400 26.200 133.000 27.600 ;
        RECT 115.800 22.200 116.600 23.600 ;
        RECT 119.600 22.200 120.400 24.200 ;
        RECT 127.600 26.000 131.600 26.200 ;
        RECT 127.600 22.200 128.400 26.000 ;
        RECT 130.800 22.200 131.600 26.000 ;
        RECT 132.400 22.200 133.200 26.200 ;
        RECT 138.400 25.000 139.000 31.600 ;
        RECT 149.800 30.400 150.600 30.600 ;
        RECT 151.800 30.400 152.400 31.800 ;
        RECT 165.000 31.600 168.400 32.200 ;
        RECT 170.800 31.800 173.000 32.400 ;
        RECT 139.600 29.600 141.200 30.400 ;
        RECT 149.000 29.800 150.600 30.400 ;
        RECT 151.600 30.300 152.400 30.400 ;
        RECT 149.000 29.600 149.800 29.800 ;
        RECT 151.600 29.700 161.900 30.300 ;
        RECT 151.600 29.600 152.400 29.700 ;
        RECT 150.400 28.600 151.200 28.800 ;
        RECT 148.400 28.400 151.200 28.600 ;
        RECT 141.200 28.300 142.800 28.400 ;
        RECT 143.600 28.300 144.400 28.400 ;
        RECT 141.200 27.700 144.400 28.300 ;
        RECT 141.200 27.600 142.800 27.700 ;
        RECT 143.600 27.600 144.400 27.700 ;
        RECT 146.800 28.000 151.200 28.400 ;
        RECT 151.800 28.400 152.400 29.600 ;
        RECT 161.300 28.400 161.900 29.700 ;
        RECT 162.800 29.600 164.400 30.400 ;
        RECT 146.800 27.800 149.000 28.000 ;
        RECT 151.800 27.800 152.800 28.400 ;
        RECT 146.800 27.600 148.400 27.800 ;
        RECT 148.600 26.800 149.400 27.000 ;
        RECT 140.400 26.300 141.200 26.400 ;
        RECT 142.600 26.300 144.400 26.400 ;
        RECT 140.400 25.700 144.400 26.300 ;
        RECT 140.400 25.600 141.200 25.700 ;
        RECT 142.600 25.600 144.400 25.700 ;
        RECT 146.800 26.200 149.400 26.800 ;
        RECT 150.000 26.400 151.600 27.200 ;
        RECT 138.400 24.400 142.400 25.000 ;
        RECT 138.400 24.200 139.600 24.400 ;
        RECT 138.800 22.200 139.600 24.200 ;
        RECT 141.800 23.600 142.800 24.400 ;
        RECT 142.000 22.200 142.800 23.600 ;
        RECT 146.800 22.200 147.600 26.200 ;
        RECT 152.200 25.800 152.800 27.800 ;
        RECT 153.600 27.600 154.400 28.400 ;
        RECT 161.200 27.600 162.800 28.400 ;
        RECT 153.600 27.200 154.200 27.600 ;
        RECT 153.400 26.400 154.200 27.200 ;
        RECT 154.800 26.800 155.600 27.000 ;
        RECT 154.800 26.200 157.200 26.800 ;
        RECT 151.200 22.200 152.800 25.800 ;
        RECT 156.400 22.200 157.200 26.200 ;
        RECT 159.600 25.600 161.400 26.400 ;
        RECT 165.000 25.000 165.600 31.600 ;
        RECT 172.400 31.200 173.000 31.800 ;
        RECT 172.400 30.400 173.600 31.200 ;
        RECT 172.400 27.400 173.000 30.400 ;
        RECT 161.600 24.400 165.600 25.000 ;
        RECT 170.800 26.800 173.000 27.400 ;
        RECT 161.600 24.200 162.200 24.400 ;
        RECT 161.200 23.600 162.200 24.200 ;
        RECT 164.400 24.300 165.600 24.400 ;
        RECT 169.200 24.300 170.000 24.400 ;
        RECT 164.400 23.700 170.000 24.300 ;
        RECT 161.200 22.200 162.000 23.600 ;
        RECT 164.400 22.200 165.200 23.700 ;
        RECT 169.200 23.600 170.000 23.700 ;
        RECT 170.800 22.200 171.600 26.800 ;
        RECT 4.400 15.200 5.200 19.800 ;
        RECT 9.200 15.200 10.000 19.800 ;
        RECT 11.400 16.800 12.200 19.800 ;
        RECT 3.000 14.600 5.200 15.200 ;
        RECT 7.800 14.600 10.000 15.200 ;
        RECT 10.800 15.800 12.200 16.800 ;
        RECT 15.600 15.800 16.400 19.800 ;
        RECT 3.000 11.600 3.600 14.600 ;
        RECT 4.400 11.600 5.200 13.200 ;
        RECT 7.800 11.600 8.400 14.600 ;
        RECT 9.200 12.300 10.000 13.200 ;
        RECT 10.800 12.400 11.400 15.800 ;
        RECT 15.600 15.600 16.200 15.800 ;
        RECT 14.400 15.200 16.200 15.600 ;
        RECT 20.400 15.200 21.200 19.800 ;
        RECT 25.200 18.400 26.000 19.800 ;
        RECT 25.200 17.600 26.200 18.400 ;
        RECT 28.400 17.800 29.200 19.800 ;
        RECT 28.400 17.600 29.600 17.800 ;
        RECT 25.600 17.000 29.600 17.600 ;
        RECT 23.600 16.300 25.400 16.400 ;
        RECT 26.800 16.300 27.600 16.400 ;
        RECT 23.600 15.700 27.600 16.300 ;
        RECT 23.600 15.600 25.400 15.700 ;
        RECT 26.800 15.600 27.600 15.700 ;
        RECT 12.000 15.000 16.200 15.200 ;
        RECT 12.000 14.600 15.000 15.000 ;
        RECT 19.000 14.600 21.200 15.200 ;
        RECT 12.000 14.400 12.800 14.600 ;
        RECT 10.800 12.300 11.600 12.400 ;
        RECT 9.200 11.700 11.600 12.300 ;
        RECT 9.200 11.600 10.000 11.700 ;
        RECT 10.800 11.600 11.600 11.700 ;
        RECT 2.400 10.800 3.600 11.600 ;
        RECT 7.200 10.800 8.400 11.600 ;
        RECT 3.000 10.200 3.600 10.800 ;
        RECT 7.800 10.200 8.400 10.800 ;
        RECT 10.800 10.200 11.400 11.600 ;
        RECT 12.200 11.000 12.800 14.400 ;
        RECT 13.600 13.800 14.400 14.000 ;
        RECT 13.600 13.200 14.600 13.800 ;
        RECT 14.000 12.400 14.600 13.200 ;
        RECT 15.600 12.800 16.400 14.400 ;
        RECT 14.000 11.600 14.800 12.400 ;
        RECT 19.000 11.600 19.600 14.600 ;
        RECT 22.000 14.300 22.800 14.400 ;
        RECT 25.200 14.300 26.800 14.400 ;
        RECT 22.000 13.700 26.800 14.300 ;
        RECT 22.000 13.600 22.800 13.700 ;
        RECT 25.200 13.600 26.800 13.700 ;
        RECT 20.400 12.300 21.200 13.200 ;
        RECT 25.200 12.300 26.000 12.400 ;
        RECT 20.400 11.700 26.000 12.300 ;
        RECT 20.400 11.600 21.200 11.700 ;
        RECT 25.200 11.600 26.000 11.700 ;
        RECT 26.800 11.600 28.400 12.400 ;
        RECT 12.200 10.400 14.600 11.000 ;
        RECT 18.400 10.800 19.600 11.600 ;
        RECT 3.000 9.600 5.200 10.200 ;
        RECT 7.800 9.600 10.000 10.200 ;
        RECT 4.400 2.200 5.200 9.600 ;
        RECT 9.200 2.200 10.000 9.600 ;
        RECT 10.800 2.200 11.600 10.200 ;
        RECT 14.000 6.200 14.600 10.400 ;
        RECT 19.000 10.200 19.600 10.800 ;
        RECT 29.000 10.400 29.600 17.000 ;
        RECT 38.000 15.200 38.800 19.800 ;
        RECT 42.800 18.400 43.600 19.800 ;
        RECT 42.800 17.600 43.800 18.400 ;
        RECT 46.000 17.800 46.800 19.800 ;
        RECT 46.000 17.600 47.200 17.800 ;
        RECT 43.200 17.000 47.200 17.600 ;
        RECT 41.200 16.300 43.000 16.400 ;
        RECT 44.400 16.300 45.200 16.400 ;
        RECT 41.200 15.700 45.200 16.300 ;
        RECT 41.200 15.600 43.000 15.700 ;
        RECT 44.400 15.600 45.200 15.700 ;
        RECT 36.600 14.600 38.800 15.200 ;
        RECT 36.600 11.600 37.200 14.600 ;
        RECT 42.800 13.600 44.400 14.400 ;
        RECT 38.000 12.300 38.800 13.200 ;
        RECT 41.200 12.300 42.000 12.400 ;
        RECT 38.000 11.700 42.000 12.300 ;
        RECT 38.000 11.600 38.800 11.700 ;
        RECT 41.200 11.600 42.000 11.700 ;
        RECT 44.400 11.600 46.000 12.400 ;
        RECT 36.000 10.800 37.200 11.600 ;
        RECT 19.000 9.600 21.200 10.200 ;
        RECT 29.000 9.800 32.400 10.400 ;
        RECT 14.000 2.200 14.800 6.200 ;
        RECT 20.400 2.200 21.200 9.600 ;
        RECT 31.600 9.600 32.400 9.800 ;
        RECT 36.600 10.200 37.200 10.800 ;
        RECT 46.600 10.400 47.200 17.000 ;
        RECT 57.200 15.200 58.000 19.800 ;
        RECT 63.600 17.800 64.400 19.800 ;
        RECT 67.400 18.400 68.200 19.800 ;
        RECT 57.200 14.600 59.400 15.200 ;
        RECT 57.200 11.600 58.000 13.200 ;
        RECT 58.800 11.600 59.400 14.600 ;
        RECT 63.600 14.400 64.200 17.800 ;
        RECT 66.800 17.600 68.200 18.400 ;
        RECT 67.400 16.800 68.200 17.600 ;
        RECT 66.800 15.800 68.200 16.800 ;
        RECT 71.600 15.800 72.400 19.800 ;
        RECT 73.800 18.400 74.600 19.800 ;
        RECT 73.200 17.600 74.600 18.400 ;
        RECT 82.800 17.800 83.600 19.800 ;
        RECT 86.000 18.400 86.800 19.800 ;
        RECT 73.800 16.400 74.600 17.600 ;
        RECT 82.400 17.600 83.600 17.800 ;
        RECT 85.800 17.600 86.800 18.400 ;
        RECT 82.400 17.000 86.400 17.600 ;
        RECT 73.800 15.800 75.600 16.400 ;
        RECT 63.600 13.600 64.400 14.400 ;
        RECT 63.600 12.400 64.200 13.600 ;
        RECT 66.800 12.400 67.400 15.800 ;
        RECT 71.600 15.600 72.200 15.800 ;
        RECT 70.400 15.200 72.200 15.600 ;
        RECT 68.000 15.000 72.200 15.200 ;
        RECT 68.000 14.600 71.000 15.000 ;
        RECT 68.000 14.400 68.800 14.600 ;
        RECT 63.600 11.600 64.400 12.400 ;
        RECT 66.800 11.600 67.600 12.400 ;
        RECT 58.800 10.800 60.000 11.600 ;
        RECT 36.600 9.600 38.800 10.200 ;
        RECT 46.600 9.800 50.000 10.400 ;
        RECT 58.800 10.200 59.400 10.800 ;
        RECT 63.600 10.200 64.200 11.600 ;
        RECT 66.800 10.200 67.400 11.600 ;
        RECT 68.200 11.000 68.800 14.400 ;
        RECT 69.600 13.800 70.400 14.000 ;
        RECT 69.600 13.200 70.600 13.800 ;
        RECT 70.000 12.400 70.600 13.200 ;
        RECT 71.600 12.800 72.400 14.400 ;
        RECT 70.000 11.600 70.800 12.400 ;
        RECT 68.200 10.400 70.600 11.000 ;
        RECT 22.200 8.800 25.800 9.400 ;
        RECT 22.200 8.200 22.800 8.800 ;
        RECT 22.000 2.200 22.800 8.200 ;
        RECT 25.200 8.200 25.800 8.800 ;
        RECT 27.000 9.000 30.600 9.200 ;
        RECT 31.600 9.000 32.200 9.600 ;
        RECT 27.000 8.600 30.800 9.000 ;
        RECT 27.000 8.200 27.600 8.600 ;
        RECT 25.200 2.800 26.000 8.200 ;
        RECT 26.800 3.400 27.600 8.200 ;
        RECT 28.400 2.800 29.200 8.000 ;
        RECT 30.000 3.000 30.800 8.600 ;
        RECT 31.600 3.400 32.400 9.000 ;
        RECT 25.200 2.200 29.200 2.800 ;
        RECT 30.200 2.800 30.800 3.000 ;
        RECT 33.200 3.000 34.000 9.000 ;
        RECT 33.200 2.800 33.800 3.000 ;
        RECT 30.200 2.200 33.800 2.800 ;
        RECT 38.000 2.200 38.800 9.600 ;
        RECT 49.200 9.600 50.000 9.800 ;
        RECT 57.200 9.600 59.400 10.200 ;
        RECT 39.800 8.800 43.400 9.400 ;
        RECT 39.800 8.200 40.400 8.800 ;
        RECT 39.600 2.200 40.400 8.200 ;
        RECT 42.800 8.200 43.400 8.800 ;
        RECT 44.600 9.000 48.200 9.200 ;
        RECT 49.200 9.000 49.800 9.600 ;
        RECT 44.600 8.600 48.400 9.000 ;
        RECT 44.600 8.200 45.200 8.600 ;
        RECT 42.800 2.800 43.600 8.200 ;
        RECT 44.400 3.400 45.200 8.200 ;
        RECT 46.000 2.800 46.800 8.000 ;
        RECT 47.600 3.000 48.400 8.600 ;
        RECT 49.200 3.400 50.000 9.000 ;
        RECT 42.800 2.200 46.800 2.800 ;
        RECT 47.800 2.800 48.400 3.000 ;
        RECT 50.800 3.000 51.600 9.000 ;
        RECT 50.800 2.800 51.400 3.000 ;
        RECT 47.800 2.200 51.400 2.800 ;
        RECT 57.200 2.200 58.000 9.600 ;
        RECT 62.600 9.400 64.400 10.200 ;
        RECT 62.600 2.200 63.400 9.400 ;
        RECT 66.800 2.200 67.600 10.200 ;
        RECT 70.000 6.200 70.600 10.400 ;
        RECT 73.200 8.800 74.000 10.400 ;
        RECT 70.000 2.200 70.800 6.200 ;
        RECT 74.800 2.200 75.600 15.800 ;
        RECT 76.400 13.600 77.200 15.200 ;
        RECT 82.400 10.400 83.000 17.000 ;
        RECT 86.600 16.300 88.400 16.400 ;
        RECT 89.200 16.300 90.000 16.400 ;
        RECT 86.600 15.700 90.000 16.300 ;
        RECT 86.600 15.600 88.400 15.700 ;
        RECT 89.200 15.600 90.000 15.700 ;
        RECT 90.800 15.200 91.600 19.800 ;
        RECT 97.200 17.600 98.000 19.800 ;
        RECT 90.800 14.600 93.000 15.200 ;
        RECT 85.200 14.300 86.800 14.400 ;
        RECT 87.600 14.300 88.400 14.400 ;
        RECT 85.200 13.700 88.400 14.300 ;
        RECT 85.200 13.600 86.800 13.700 ;
        RECT 87.600 13.600 88.400 13.700 ;
        RECT 83.600 11.600 85.200 12.400 ;
        RECT 86.000 12.300 86.800 12.400 ;
        RECT 90.800 12.300 91.600 13.200 ;
        RECT 86.000 11.700 91.600 12.300 ;
        RECT 86.000 11.600 86.800 11.700 ;
        RECT 90.800 11.600 91.600 11.700 ;
        RECT 92.400 11.600 93.000 14.600 ;
        RECT 97.400 14.400 98.000 17.600 ;
        RECT 100.400 15.800 101.200 19.800 ;
        RECT 104.800 18.400 106.400 19.800 ;
        RECT 104.800 17.600 107.600 18.400 ;
        RECT 104.800 16.200 106.400 17.600 ;
        RECT 100.400 15.200 102.800 15.800 ;
        RECT 102.000 15.000 102.800 15.200 ;
        RECT 103.400 14.800 104.200 15.600 ;
        RECT 103.400 14.400 104.000 14.800 ;
        RECT 97.200 13.600 98.000 14.400 ;
        RECT 103.200 13.600 104.000 14.400 ;
        RECT 104.800 14.200 105.400 16.200 ;
        RECT 110.000 15.800 110.800 19.800 ;
        RECT 106.000 14.800 107.600 15.600 ;
        RECT 108.200 15.200 110.800 15.800 ;
        RECT 111.600 15.800 112.400 19.800 ;
        RECT 116.000 16.200 117.600 19.800 ;
        RECT 111.600 15.200 114.200 15.800 ;
        RECT 108.200 15.000 109.000 15.200 ;
        RECT 113.400 15.000 114.200 15.200 ;
        RECT 114.800 14.800 116.400 15.600 ;
        RECT 109.200 14.200 110.800 14.400 ;
        RECT 104.800 13.600 105.800 14.200 ;
        RECT 108.600 14.000 110.800 14.200 ;
        RECT 79.600 9.800 83.000 10.400 ;
        RECT 92.400 10.800 93.600 11.600 ;
        RECT 92.400 10.200 93.000 10.800 ;
        RECT 97.400 10.200 98.000 13.600 ;
        RECT 105.200 12.400 105.800 13.600 ;
        RECT 106.400 13.600 110.800 14.000 ;
        RECT 111.600 14.200 113.200 14.400 ;
        RECT 117.000 14.200 117.600 16.200 ;
        RECT 121.200 15.800 122.000 19.800 ;
        RECT 132.400 17.800 133.200 19.800 ;
        RECT 135.600 18.400 136.400 19.800 ;
        RECT 118.200 14.800 119.000 15.600 ;
        RECT 119.600 15.200 122.000 15.800 ;
        RECT 132.000 17.600 133.200 17.800 ;
        RECT 135.400 17.800 136.400 18.400 ;
        RECT 135.400 17.600 136.000 17.800 ;
        RECT 132.000 17.000 136.000 17.600 ;
        RECT 119.600 15.000 120.400 15.200 ;
        RECT 111.600 14.000 113.800 14.200 ;
        RECT 111.600 13.600 116.000 14.000 ;
        RECT 106.400 13.400 109.200 13.600 ;
        RECT 113.200 13.400 116.000 13.600 ;
        RECT 106.400 13.200 107.200 13.400 ;
        RECT 115.200 13.200 116.000 13.400 ;
        RECT 116.600 13.600 117.600 14.200 ;
        RECT 118.400 14.400 119.000 14.800 ;
        RECT 132.000 14.400 132.600 17.000 ;
        RECT 135.600 15.600 138.000 16.400 ;
        RECT 140.400 15.200 141.200 19.800 ;
        RECT 145.200 15.200 146.000 19.800 ;
        RECT 154.800 17.800 155.600 19.800 ;
        RECT 158.000 18.400 158.800 19.800 ;
        RECT 154.400 17.600 155.600 17.800 ;
        RECT 157.800 17.800 158.800 18.400 ;
        RECT 157.800 17.600 158.400 17.800 ;
        RECT 154.400 17.000 158.400 17.600 ;
        RECT 140.400 14.600 142.600 15.200 ;
        RECT 145.200 14.600 147.400 15.200 ;
        RECT 118.400 13.600 119.200 14.400 ;
        RECT 132.000 13.600 133.200 14.400 ;
        RECT 134.800 13.600 136.400 14.400 ;
        RECT 116.600 12.400 117.200 13.600 ;
        RECT 105.200 11.600 106.000 12.400 ;
        RECT 107.800 12.200 108.600 12.400 ;
        RECT 107.000 11.600 108.600 12.200 ;
        RECT 113.800 12.200 114.600 12.400 ;
        RECT 116.400 12.300 117.200 12.400 ;
        RECT 129.200 12.300 130.000 12.400 ;
        RECT 113.800 11.600 115.400 12.200 ;
        RECT 116.400 11.700 130.000 12.300 ;
        RECT 116.400 11.600 117.200 11.700 ;
        RECT 129.200 11.600 130.000 11.700 ;
        RECT 105.200 10.200 105.800 11.600 ;
        RECT 107.000 11.400 107.800 11.600 ;
        RECT 114.600 11.400 115.400 11.600 ;
        RECT 116.600 10.200 117.200 11.600 ;
        RECT 132.000 10.400 132.600 13.600 ;
        RECT 133.200 11.600 134.800 12.400 ;
        RECT 140.400 11.600 141.200 13.200 ;
        RECT 142.000 11.600 142.600 14.600 ;
        RECT 145.200 11.600 146.000 13.200 ;
        RECT 146.800 11.600 147.400 14.600 ;
        RECT 154.400 14.400 155.000 17.000 ;
        RECT 158.000 15.600 160.400 16.400 ;
        RECT 162.800 15.200 163.600 19.800 ;
        RECT 168.200 18.400 169.000 19.800 ;
        RECT 167.600 17.600 169.000 18.400 ;
        RECT 168.200 16.800 169.000 17.600 ;
        RECT 167.600 15.800 169.000 16.800 ;
        RECT 172.400 15.800 173.200 19.800 ;
        RECT 162.800 14.600 165.000 15.200 ;
        RECT 154.400 13.600 155.600 14.400 ;
        RECT 157.200 14.300 158.800 14.400 ;
        RECT 159.600 14.300 160.400 14.400 ;
        RECT 157.200 13.700 160.400 14.300 ;
        RECT 157.200 13.600 158.800 13.700 ;
        RECT 159.600 13.600 160.400 13.700 ;
        RECT 79.600 9.600 80.400 9.800 ;
        RECT 79.800 9.000 80.400 9.600 ;
        RECT 90.800 9.600 93.000 10.200 ;
        RECT 81.400 9.000 85.000 9.200 ;
        RECT 78.000 3.000 78.800 9.000 ;
        RECT 79.600 3.400 80.400 9.000 ;
        RECT 81.200 8.600 85.000 9.000 ;
        RECT 78.200 2.800 78.800 3.000 ;
        RECT 81.200 3.000 82.000 8.600 ;
        RECT 84.400 8.200 85.000 8.600 ;
        RECT 86.200 8.800 89.800 9.400 ;
        RECT 86.200 8.200 86.800 8.800 ;
        RECT 81.200 2.800 81.800 3.000 ;
        RECT 78.200 2.200 81.800 2.800 ;
        RECT 82.800 2.800 83.600 8.000 ;
        RECT 84.400 3.400 85.200 8.200 ;
        RECT 86.000 2.800 86.800 8.200 ;
        RECT 82.800 2.200 86.800 2.800 ;
        RECT 89.200 8.200 89.800 8.800 ;
        RECT 89.200 2.200 90.000 8.200 ;
        RECT 90.800 2.200 91.600 9.600 ;
        RECT 97.200 9.400 99.000 10.200 ;
        RECT 98.200 2.200 99.000 9.400 ;
        RECT 100.400 9.600 102.800 10.200 ;
        RECT 100.400 2.200 101.200 9.600 ;
        RECT 102.000 9.400 102.800 9.600 ;
        RECT 104.800 2.200 106.400 10.200 ;
        RECT 108.200 9.600 110.800 10.200 ;
        RECT 108.200 9.400 109.000 9.600 ;
        RECT 110.000 2.200 110.800 9.600 ;
        RECT 111.600 9.600 114.200 10.200 ;
        RECT 111.600 2.200 112.400 9.600 ;
        RECT 113.400 9.400 114.200 9.600 ;
        RECT 116.000 2.200 117.600 10.200 ;
        RECT 119.600 9.600 122.000 10.200 ;
        RECT 129.200 9.800 132.600 10.400 ;
        RECT 142.000 10.800 143.200 11.600 ;
        RECT 146.800 10.800 148.000 11.600 ;
        RECT 142.000 10.200 142.600 10.800 ;
        RECT 146.800 10.200 147.400 10.800 ;
        RECT 154.400 10.400 155.000 13.600 ;
        RECT 155.600 12.300 157.200 12.400 ;
        RECT 161.200 12.300 162.000 12.400 ;
        RECT 155.600 11.700 162.000 12.300 ;
        RECT 155.600 11.600 157.200 11.700 ;
        RECT 161.200 11.600 162.000 11.700 ;
        RECT 162.800 11.600 163.600 13.200 ;
        RECT 164.400 11.600 165.000 14.600 ;
        RECT 167.600 12.400 168.200 15.800 ;
        RECT 172.400 15.600 173.000 15.800 ;
        RECT 171.200 15.200 173.000 15.600 ;
        RECT 177.200 15.200 178.000 19.800 ;
        RECT 168.800 15.000 173.000 15.200 ;
        RECT 168.800 14.600 171.800 15.000 ;
        RECT 175.800 14.600 178.000 15.200 ;
        RECT 168.800 14.400 169.600 14.600 ;
        RECT 167.600 11.600 168.400 12.400 ;
        RECT 129.200 9.600 130.000 9.800 ;
        RECT 119.600 9.400 120.400 9.600 ;
        RECT 121.200 2.200 122.000 9.600 ;
        RECT 129.400 9.000 130.000 9.600 ;
        RECT 140.400 9.600 142.600 10.200 ;
        RECT 145.200 9.600 147.400 10.200 ;
        RECT 151.600 9.800 155.000 10.400 ;
        RECT 164.400 10.800 165.600 11.600 ;
        RECT 164.400 10.200 165.000 10.800 ;
        RECT 151.600 9.600 152.400 9.800 ;
        RECT 131.000 9.000 134.600 9.200 ;
        RECT 127.600 3.000 128.400 9.000 ;
        RECT 129.200 3.400 130.000 9.000 ;
        RECT 130.800 8.600 134.600 9.000 ;
        RECT 127.800 2.800 128.400 3.000 ;
        RECT 130.800 3.000 131.600 8.600 ;
        RECT 134.000 8.200 134.600 8.600 ;
        RECT 135.800 8.800 139.400 9.400 ;
        RECT 135.800 8.200 136.400 8.800 ;
        RECT 130.800 2.800 131.400 3.000 ;
        RECT 127.800 2.200 131.400 2.800 ;
        RECT 132.400 2.800 133.200 8.000 ;
        RECT 134.000 3.400 134.800 8.200 ;
        RECT 135.600 2.800 136.400 8.200 ;
        RECT 132.400 2.200 136.400 2.800 ;
        RECT 138.800 8.200 139.400 8.800 ;
        RECT 138.800 2.200 139.600 8.200 ;
        RECT 140.400 2.200 141.200 9.600 ;
        RECT 145.200 2.200 146.000 9.600 ;
        RECT 151.800 9.000 152.400 9.600 ;
        RECT 162.800 9.600 165.000 10.200 ;
        RECT 167.600 10.200 168.200 11.600 ;
        RECT 169.000 11.000 169.600 14.400 ;
        RECT 170.400 13.800 171.200 14.000 ;
        RECT 170.400 13.200 171.400 13.800 ;
        RECT 170.800 12.400 171.400 13.200 ;
        RECT 172.400 12.800 173.200 14.400 ;
        RECT 170.800 11.600 171.600 12.400 ;
        RECT 175.800 11.600 176.400 14.600 ;
        RECT 177.200 11.600 178.000 13.200 ;
        RECT 169.000 10.400 171.400 11.000 ;
        RECT 175.200 10.800 176.400 11.600 ;
        RECT 153.400 9.000 157.000 9.200 ;
        RECT 150.000 3.000 150.800 9.000 ;
        RECT 151.600 3.400 152.400 9.000 ;
        RECT 153.200 8.600 157.000 9.000 ;
        RECT 150.200 2.800 150.800 3.000 ;
        RECT 153.200 3.000 154.000 8.600 ;
        RECT 156.400 8.200 157.000 8.600 ;
        RECT 158.200 8.800 161.800 9.400 ;
        RECT 158.200 8.200 158.800 8.800 ;
        RECT 153.200 2.800 153.800 3.000 ;
        RECT 150.200 2.200 153.800 2.800 ;
        RECT 154.800 2.800 155.600 8.000 ;
        RECT 156.400 3.400 157.200 8.200 ;
        RECT 158.000 2.800 158.800 8.200 ;
        RECT 154.800 2.200 158.800 2.800 ;
        RECT 161.200 8.200 161.800 8.800 ;
        RECT 161.200 2.200 162.000 8.200 ;
        RECT 162.800 2.200 163.600 9.600 ;
        RECT 167.600 2.200 168.400 10.200 ;
        RECT 170.800 6.200 171.400 10.400 ;
        RECT 175.800 10.200 176.400 10.800 ;
        RECT 175.800 9.600 178.000 10.200 ;
        RECT 170.800 2.200 171.600 6.200 ;
        RECT 177.200 2.200 178.000 9.600 ;
      LAYER via1 ;
        RECT 10.800 133.600 11.600 134.400 ;
        RECT 6.000 123.600 6.800 124.400 ;
        RECT 60.400 133.600 61.200 134.400 ;
        RECT 63.600 133.600 64.400 134.400 ;
        RECT 49.200 131.600 50.000 132.400 ;
        RECT 62.000 131.600 62.800 132.400 ;
        RECT 74.800 133.600 75.600 134.400 ;
        RECT 84.400 133.600 85.200 134.400 ;
        RECT 73.200 131.600 74.000 132.400 ;
        RECT 76.400 131.600 77.200 132.400 ;
        RECT 87.600 133.600 88.400 134.400 ;
        RECT 81.200 123.600 82.000 124.400 ;
        RECT 98.800 134.800 99.600 135.600 ;
        RECT 102.000 131.600 102.800 132.400 ;
        RECT 124.400 135.600 125.200 136.400 ;
        RECT 119.600 133.600 120.400 134.400 ;
        RECT 122.800 133.600 123.600 134.400 ;
        RECT 121.200 131.600 122.000 132.400 ;
        RECT 111.600 123.600 112.400 124.400 ;
        RECT 1.200 107.600 2.000 108.400 ;
        RECT 28.400 111.800 29.200 112.600 ;
        RECT 17.200 109.600 18.000 110.400 ;
        RECT 12.400 107.600 13.200 108.400 ;
        RECT 15.600 107.600 16.400 108.400 ;
        RECT 4.400 103.600 5.200 104.400 ;
        RECT 10.800 105.600 11.600 106.400 ;
        RECT 18.800 107.600 19.600 108.400 ;
        RECT 28.400 106.200 29.200 107.000 ;
        RECT 25.200 103.600 26.000 104.400 ;
        RECT 33.200 106.400 34.000 107.200 ;
        RECT 33.200 103.600 34.000 104.400 ;
        RECT 42.800 105.600 43.600 106.400 ;
        RECT 70.000 111.600 70.800 112.400 ;
        RECT 65.200 109.600 66.000 110.400 ;
        RECT 57.200 107.600 58.000 108.400 ;
        RECT 58.800 107.600 59.600 108.400 ;
        RECT 66.800 107.600 67.600 108.400 ;
        RECT 71.600 107.600 72.400 108.400 ;
        RECT 54.000 103.600 54.800 104.400 ;
        RECT 101.800 111.800 102.600 112.600 ;
        RECT 113.200 117.600 114.000 118.400 ;
        RECT 130.800 117.600 131.600 118.400 ;
        RECT 95.600 109.600 96.400 110.400 ;
        RECT 79.600 105.600 80.400 106.400 ;
        RECT 101.800 106.200 102.600 107.000 ;
        RECT 119.600 107.600 120.400 108.400 ;
        RECT 135.600 109.600 136.400 110.400 ;
        RECT 137.200 107.600 138.000 108.400 ;
        RECT 148.400 109.600 149.200 110.400 ;
        RECT 150.000 107.600 150.800 108.400 ;
        RECT 158.000 107.600 158.800 108.400 ;
        RECT 166.000 109.600 166.800 110.400 ;
        RECT 31.600 94.800 32.400 95.600 ;
        RECT 15.600 89.600 16.400 90.400 ;
        RECT 26.800 89.600 27.600 90.400 ;
        RECT 34.800 89.600 35.600 90.400 ;
        RECT 62.000 89.600 62.800 90.400 ;
        RECT 57.200 83.600 58.000 84.400 ;
        RECT 63.600 89.600 64.400 90.400 ;
        RECT 95.600 95.600 96.400 96.400 ;
        RECT 78.000 91.600 78.800 92.400 ;
        RECT 66.800 83.600 67.600 84.400 ;
        RECT 87.600 91.600 88.400 92.400 ;
        RECT 119.600 97.600 120.400 98.400 ;
        RECT 114.800 91.600 115.600 92.400 ;
        RECT 137.200 97.600 138.000 98.400 ;
        RECT 114.800 83.600 115.600 84.400 ;
        RECT 143.600 93.600 144.400 94.400 ;
        RECT 124.400 89.600 125.200 90.400 ;
        RECT 148.400 89.600 149.200 90.400 ;
        RECT 154.800 83.600 155.600 84.400 ;
        RECT 161.200 89.600 162.000 90.400 ;
        RECT 159.600 83.600 160.400 84.400 ;
        RECT 7.600 73.600 8.400 74.400 ;
        RECT 18.800 77.600 19.600 78.400 ;
        RECT 23.600 77.600 24.400 78.400 ;
        RECT 17.200 73.600 18.000 74.400 ;
        RECT 25.200 73.600 26.000 74.400 ;
        RECT 30.000 73.600 30.800 74.400 ;
        RECT 20.400 71.600 21.200 72.400 ;
        RECT 22.000 71.600 22.800 72.400 ;
        RECT 18.800 69.600 19.600 70.400 ;
        RECT 9.200 65.600 10.000 66.400 ;
        RECT 33.200 71.600 34.000 72.400 ;
        RECT 36.400 71.800 37.200 72.600 ;
        RECT 31.600 69.600 32.400 70.400 ;
        RECT 36.400 66.200 37.200 67.000 ;
        RECT 54.000 69.600 54.800 70.400 ;
        RECT 70.000 73.600 70.800 74.400 ;
        RECT 66.800 71.600 67.600 72.400 ;
        RECT 65.200 69.600 66.000 70.400 ;
        RECT 41.200 66.400 42.000 67.200 ;
        RECT 41.200 63.600 42.000 64.400 ;
        RECT 82.800 75.600 83.600 76.400 ;
        RECT 92.400 77.600 93.200 78.400 ;
        RECT 89.200 73.600 90.000 74.400 ;
        RECT 86.000 71.600 86.800 72.400 ;
        RECT 76.400 67.600 77.200 68.400 ;
        RECT 97.200 71.800 98.000 72.600 ;
        RECT 113.200 77.600 114.000 78.400 ;
        RECT 121.200 77.600 122.000 78.400 ;
        RECT 110.000 69.600 110.800 70.400 ;
        RECT 94.000 65.600 94.800 66.400 ;
        RECT 97.200 66.200 98.000 67.000 ;
        RECT 92.400 63.600 93.200 64.400 ;
        RECT 102.000 66.400 102.800 67.200 ;
        RECT 111.600 67.600 112.400 68.400 ;
        RECT 113.200 63.600 114.000 64.400 ;
        RECT 121.200 63.600 122.000 64.400 ;
        RECT 132.400 67.600 133.200 68.400 ;
        RECT 137.200 67.600 138.000 68.400 ;
        RECT 150.200 71.800 151.000 72.600 ;
        RECT 162.800 77.600 163.600 78.400 ;
        RECT 145.200 69.600 146.000 70.400 ;
        RECT 151.400 69.800 152.200 70.600 ;
        RECT 143.600 67.600 144.400 68.400 ;
        RECT 150.200 66.200 151.000 67.000 ;
        RECT 140.400 63.600 141.200 64.400 ;
        RECT 154.800 63.600 155.600 64.400 ;
        RECT 161.200 63.600 162.000 64.400 ;
        RECT 12.400 57.600 13.200 58.400 ;
        RECT 20.400 57.600 21.200 58.400 ;
        RECT 10.800 49.600 11.600 50.400 ;
        RECT 15.600 53.600 16.400 54.400 ;
        RECT 28.400 54.800 29.200 55.600 ;
        RECT 31.600 53.600 32.400 54.400 ;
        RECT 41.200 53.600 42.000 54.400 ;
        RECT 39.600 51.600 40.400 52.400 ;
        RECT 42.800 51.600 43.600 52.400 ;
        RECT 68.400 57.600 69.200 58.400 ;
        RECT 54.000 45.600 54.800 46.400 ;
        RECT 63.600 49.600 64.400 50.400 ;
        RECT 68.400 49.600 69.200 50.400 ;
        RECT 84.400 57.600 85.200 58.400 ;
        RECT 95.600 57.600 96.400 58.400 ;
        RECT 73.200 51.600 74.000 52.400 ;
        RECT 70.000 43.600 70.800 44.400 ;
        RECT 78.000 43.600 78.800 44.400 ;
        RECT 82.800 49.600 83.600 50.400 ;
        RECT 97.200 55.600 98.000 56.400 ;
        RECT 100.400 49.600 101.200 50.400 ;
        RECT 102.000 43.600 102.800 44.400 ;
        RECT 110.000 53.600 110.800 54.400 ;
        RECT 111.600 49.600 112.400 50.400 ;
        RECT 116.400 49.600 117.200 50.400 ;
        RECT 118.000 43.600 118.800 44.400 ;
        RECT 134.000 53.600 134.800 54.400 ;
        RECT 135.600 51.600 136.400 52.400 ;
        RECT 121.200 47.600 122.000 48.400 ;
        RECT 7.600 29.600 8.400 30.400 ;
        RECT 9.200 27.600 10.000 28.400 ;
        RECT 10.800 25.600 11.600 26.400 ;
        RECT 22.000 29.600 22.800 30.400 ;
        RECT 17.200 27.600 18.000 28.400 ;
        RECT 14.000 23.600 14.800 24.400 ;
        RECT 31.600 33.600 32.400 34.400 ;
        RECT 34.800 31.600 35.600 32.400 ;
        RECT 44.200 31.800 45.000 32.600 ;
        RECT 26.800 25.600 27.600 26.400 ;
        RECT 44.200 26.200 45.000 27.000 ;
        RECT 65.200 29.600 66.000 30.400 ;
        RECT 82.800 31.800 83.600 32.600 ;
        RECT 68.400 25.600 69.200 26.400 ;
        RECT 76.400 29.600 77.200 30.400 ;
        RECT 82.800 26.200 83.600 27.000 ;
        RECT 90.800 27.600 91.600 28.400 ;
        RECT 87.600 26.400 88.400 27.200 ;
        RECT 95.600 29.600 96.400 30.400 ;
        RECT 102.000 29.600 102.800 30.400 ;
        RECT 103.600 29.600 104.400 30.400 ;
        RECT 87.600 23.600 88.400 24.400 ;
        RECT 97.200 25.600 98.000 26.400 ;
        RECT 110.000 27.600 110.800 28.400 ;
        RECT 113.200 27.600 114.000 28.400 ;
        RECT 129.200 29.600 130.000 30.400 ;
        RECT 148.600 31.800 149.400 32.600 ;
        RECT 140.400 29.600 141.200 30.400 ;
        RECT 149.800 29.800 150.600 30.600 ;
        RECT 148.600 26.200 149.400 27.000 ;
        RECT 142.000 23.600 142.800 24.400 ;
        RECT 15.600 13.600 16.400 14.400 ;
        RECT 86.000 17.600 86.800 18.400 ;
        RECT 71.600 13.600 72.400 14.400 ;
        RECT 73.200 9.600 74.000 10.400 ;
        RECT 84.400 11.600 85.200 12.400 ;
        RECT 106.800 17.600 107.600 18.400 ;
        RECT 106.800 14.800 107.600 15.600 ;
        RECT 110.000 13.600 110.800 14.400 ;
        RECT 132.400 13.600 133.200 14.400 ;
        RECT 135.600 13.600 136.400 14.400 ;
        RECT 134.000 11.600 134.800 12.400 ;
        RECT 154.800 13.600 155.600 14.400 ;
        RECT 172.400 13.600 173.200 14.400 ;
      LAYER metal2 ;
        RECT 74.800 137.600 75.600 138.400 ;
        RECT 20.400 135.600 21.200 136.400 ;
        RECT 28.400 135.600 29.200 136.400 ;
        RECT 30.000 135.600 30.800 136.400 ;
        RECT 49.200 135.600 50.000 136.400 ;
        RECT 62.000 135.600 62.800 136.400 ;
        RECT 10.800 133.600 11.600 134.400 ;
        RECT 9.200 131.600 10.000 132.400 ;
        RECT 10.900 128.400 11.500 133.600 ;
        RECT 28.500 132.400 29.100 135.600 ;
        RECT 49.300 132.400 49.900 135.600 ;
        RECT 57.200 133.600 58.000 134.400 ;
        RECT 60.400 133.600 61.200 134.400 ;
        RECT 62.100 134.300 62.700 135.600 ;
        RECT 74.900 134.400 75.500 137.600 ;
        RECT 97.000 135.000 97.800 135.800 ;
        RECT 98.800 135.000 103.000 135.600 ;
        RECT 103.600 135.000 104.400 135.800 ;
        RECT 124.400 135.600 125.200 136.400 ;
        RECT 63.600 134.300 64.400 134.400 ;
        RECT 62.100 133.700 64.400 134.300 ;
        RECT 63.600 133.600 64.400 133.700 ;
        RECT 74.800 133.600 75.600 134.400 ;
        RECT 78.000 133.600 78.800 134.400 ;
        RECT 82.800 133.600 83.600 134.400 ;
        RECT 84.400 133.600 85.200 134.400 ;
        RECT 87.600 133.600 88.400 134.400 ;
        RECT 90.800 133.600 91.600 134.400 ;
        RECT 95.600 133.600 96.400 134.400 ;
        RECT 12.400 131.600 13.200 132.400 ;
        RECT 17.200 131.600 18.000 132.400 ;
        RECT 28.400 131.600 29.200 132.400 ;
        RECT 33.200 131.600 34.000 132.400 ;
        RECT 34.800 131.600 35.600 132.400 ;
        RECT 49.200 131.600 50.000 132.400 ;
        RECT 23.600 129.600 24.400 130.400 ;
        RECT 28.500 128.400 29.100 131.600 ;
        RECT 34.900 130.400 35.500 131.600 ;
        RECT 34.800 129.600 35.600 130.400 ;
        RECT 10.800 127.600 11.600 128.400 ;
        RECT 28.400 127.600 29.200 128.400 ;
        RECT 38.000 127.600 38.800 128.400 ;
        RECT 6.000 123.600 6.800 124.400 ;
        RECT 34.800 123.600 35.600 124.400 ;
        RECT 6.100 116.300 6.700 123.600 ;
        RECT 6.100 115.700 8.300 116.300 ;
        RECT 6.000 113.600 6.800 114.400 ;
        RECT 6.100 112.400 6.700 113.600 ;
        RECT 4.400 112.300 5.200 112.400 ;
        RECT 6.000 112.300 6.800 112.400 ;
        RECT 4.400 111.700 6.800 112.300 ;
        RECT 4.400 111.600 5.200 111.700 ;
        RECT 6.000 111.600 6.800 111.700 ;
        RECT 1.200 108.300 2.000 108.400 ;
        RECT 1.200 107.700 3.500 108.300 ;
        RECT 1.200 107.600 2.000 107.700 ;
        RECT 2.900 106.400 3.500 107.700 ;
        RECT 2.800 105.600 3.600 106.400 ;
        RECT 2.900 98.400 3.500 105.600 ;
        RECT 4.400 103.600 5.200 104.400 ;
        RECT 2.800 97.600 3.600 98.400 ;
        RECT 4.500 96.400 5.100 103.600 ;
        RECT 4.400 95.600 5.200 96.400 ;
        RECT 7.700 94.400 8.300 115.700 ;
        RECT 34.900 114.400 35.500 123.600 ;
        RECT 34.800 113.600 35.600 114.400 ;
        RECT 22.000 111.600 22.800 112.400 ;
        RECT 28.400 111.800 29.200 112.600 ;
        RECT 35.000 111.800 35.800 112.600 ;
        RECT 22.100 110.400 22.700 111.600 ;
        RECT 17.200 109.600 18.000 110.400 ;
        RECT 22.000 109.600 22.800 110.400 ;
        RECT 12.400 107.600 13.200 108.400 ;
        RECT 15.600 107.600 16.400 108.400 ;
        RECT 15.700 106.400 16.300 107.600 ;
        RECT 10.800 105.600 11.600 106.400 ;
        RECT 15.600 105.600 16.400 106.400 ;
        RECT 7.600 93.600 8.400 94.400 ;
        RECT 17.300 92.400 17.900 109.600 ;
        RECT 28.400 108.400 29.000 111.800 ;
        RECT 32.400 108.400 33.200 108.600 ;
        RECT 18.800 107.600 19.600 108.400 ;
        RECT 20.400 107.600 21.200 108.400 ;
        RECT 28.400 107.800 33.200 108.400 ;
        RECT 20.500 104.400 21.100 107.600 ;
        RECT 28.400 107.000 29.000 107.800 ;
        RECT 29.800 107.000 30.600 107.200 ;
        RECT 33.200 107.000 34.000 107.200 ;
        RECT 35.200 107.000 35.800 111.800 ;
        RECT 38.100 110.400 38.700 127.600 ;
        RECT 42.800 113.600 43.600 114.400 ;
        RECT 38.000 109.600 38.800 110.400 ;
        RECT 38.100 108.400 38.700 109.600 ;
        RECT 42.900 108.400 43.500 113.600 ;
        RECT 44.400 109.600 45.200 110.400 ;
        RECT 50.800 109.600 51.600 110.400 ;
        RECT 52.400 109.600 53.200 110.400 ;
        RECT 44.500 108.400 45.100 109.600 ;
        RECT 38.000 107.600 38.800 108.400 ;
        RECT 39.600 107.600 40.400 108.400 ;
        RECT 42.800 107.600 43.600 108.400 ;
        RECT 44.400 107.600 45.200 108.400 ;
        RECT 28.400 106.200 29.200 107.000 ;
        RECT 29.800 106.400 34.000 107.000 ;
        RECT 35.000 106.200 35.800 107.000 ;
        RECT 18.800 103.600 19.600 104.400 ;
        RECT 20.400 103.600 21.200 104.400 ;
        RECT 25.200 103.600 26.000 104.400 ;
        RECT 33.200 103.600 34.000 104.400 ;
        RECT 18.900 92.400 19.500 103.600 ;
        RECT 25.300 102.400 25.900 103.600 ;
        RECT 25.200 101.600 26.000 102.400 ;
        RECT 33.300 98.400 33.900 103.600 ;
        RECT 33.200 97.600 34.000 98.400 ;
        RECT 29.800 95.000 30.600 95.800 ;
        RECT 31.600 95.000 35.800 95.600 ;
        RECT 36.400 95.000 37.200 95.800 ;
        RECT 22.000 93.600 22.800 94.400 ;
        RECT 25.200 93.600 26.000 94.400 ;
        RECT 28.400 93.600 29.200 94.400 ;
        RECT 17.200 91.600 18.000 92.400 ;
        RECT 18.800 91.600 19.600 92.400 ;
        RECT 20.400 91.600 21.200 92.400 ;
        RECT 23.600 91.600 24.400 92.400 ;
        RECT 23.700 90.400 24.300 91.600 ;
        RECT 15.600 89.600 16.400 90.400 ;
        RECT 23.600 89.600 24.400 90.400 ;
        RECT 18.800 87.600 19.600 88.400 ;
        RECT 25.300 88.300 25.900 93.600 ;
        RECT 28.400 91.600 29.200 92.400 ;
        RECT 26.800 89.600 27.600 90.400 ;
        RECT 23.700 87.700 25.900 88.300 ;
        RECT 18.900 78.400 19.500 87.600 ;
        RECT 22.000 81.600 22.800 82.400 ;
        RECT 18.800 77.600 19.600 78.400 ;
        RECT 7.600 73.600 8.400 74.400 ;
        RECT 17.200 73.600 18.000 74.400 ;
        RECT 18.800 73.600 19.600 74.400 ;
        RECT 6.000 71.600 6.800 72.400 ;
        RECT 6.100 70.400 6.700 71.600 ;
        RECT 18.900 70.400 19.500 73.600 ;
        RECT 22.100 72.400 22.700 81.600 ;
        RECT 23.700 78.400 24.300 87.700 ;
        RECT 23.600 77.600 24.400 78.400 ;
        RECT 25.200 73.600 26.000 74.400 ;
        RECT 20.400 71.600 21.200 72.400 ;
        RECT 22.000 71.600 22.800 72.400 ;
        RECT 6.000 69.600 6.800 70.400 ;
        RECT 18.800 69.600 19.600 70.400 ;
        RECT 9.200 65.600 10.000 66.400 ;
        RECT 10.800 65.600 11.600 66.400 ;
        RECT 9.300 64.400 9.900 65.600 ;
        RECT 9.200 63.600 10.000 64.400 ;
        RECT 10.900 52.400 11.500 65.600 ;
        RECT 12.400 63.600 13.200 64.400 ;
        RECT 12.500 58.400 13.100 63.600 ;
        RECT 20.500 62.400 21.100 71.600 ;
        RECT 20.400 61.600 21.200 62.400 ;
        RECT 22.100 60.300 22.700 71.600 ;
        RECT 23.600 69.600 24.400 70.400 ;
        RECT 23.700 62.400 24.300 69.600 ;
        RECT 26.900 68.400 27.500 89.600 ;
        RECT 28.500 84.400 29.100 91.600 ;
        RECT 29.800 90.200 30.400 95.000 ;
        RECT 31.600 94.800 32.400 95.000 ;
        RECT 35.000 94.800 35.800 95.000 ;
        RECT 36.600 94.200 37.200 95.000 ;
        RECT 32.400 93.600 37.200 94.200 ;
        RECT 32.400 93.400 33.200 93.600 ;
        RECT 29.800 89.400 30.600 90.200 ;
        RECT 34.800 89.600 35.600 90.400 ;
        RECT 36.600 90.200 37.200 93.600 ;
        RECT 36.400 89.400 37.200 90.200 ;
        RECT 38.100 88.400 38.700 107.600 ;
        RECT 39.700 106.400 40.300 107.600 ;
        RECT 50.900 106.400 51.500 109.600 ;
        RECT 52.500 108.400 53.100 109.600 ;
        RECT 57.300 108.400 57.900 133.600 ;
        RECT 60.500 132.400 61.100 133.600 ;
        RECT 82.900 132.400 83.500 133.600 ;
        RECT 60.400 131.600 61.200 132.400 ;
        RECT 62.000 131.600 62.800 132.400 ;
        RECT 73.200 131.600 74.000 132.400 ;
        RECT 76.400 131.600 77.200 132.400 ;
        RECT 79.600 131.600 80.400 132.400 ;
        RECT 82.800 131.600 83.600 132.400 ;
        RECT 62.100 128.400 62.700 131.600 ;
        RECT 73.300 130.400 73.900 131.600 ;
        RECT 79.700 130.400 80.300 131.600 ;
        RECT 73.200 129.600 74.000 130.400 ;
        RECT 79.600 129.600 80.400 130.400 ;
        RECT 84.500 128.400 85.100 133.600 ;
        RECT 86.000 131.600 86.800 132.400 ;
        RECT 62.000 127.600 62.800 128.400 ;
        RECT 68.400 127.600 69.200 128.400 ;
        RECT 84.400 127.600 85.200 128.400 ;
        RECT 60.400 113.600 61.200 114.400 ;
        RECT 60.500 112.400 61.100 113.600 ;
        RECT 68.500 112.400 69.100 127.600 ;
        RECT 81.200 123.600 82.000 124.400 ;
        RECT 60.400 111.600 61.200 112.400 ;
        RECT 62.000 111.600 62.800 112.400 ;
        RECT 68.400 111.600 69.200 112.400 ;
        RECT 70.000 111.600 70.800 112.400 ;
        RECT 60.400 109.600 61.200 110.400 ;
        RECT 65.200 109.600 66.000 110.400 ;
        RECT 65.300 108.400 65.900 109.600 ;
        RECT 52.400 107.600 53.200 108.400 ;
        RECT 57.200 107.600 58.000 108.400 ;
        RECT 58.800 107.600 59.600 108.400 ;
        RECT 65.200 107.600 66.000 108.400 ;
        RECT 66.800 108.300 67.600 108.400 ;
        RECT 68.500 108.300 69.100 111.600 ;
        RECT 76.400 109.600 77.200 110.400 ;
        RECT 79.600 109.600 80.400 110.400 ;
        RECT 66.800 107.700 69.100 108.300 ;
        RECT 66.800 107.600 67.600 107.700 ;
        RECT 71.600 107.600 72.400 108.400 ;
        RECT 78.000 107.600 78.800 108.400 ;
        RECT 39.600 105.600 40.400 106.400 ;
        RECT 42.800 105.600 43.600 106.400 ;
        RECT 50.800 105.600 51.600 106.400 ;
        RECT 55.600 105.600 56.400 106.400 ;
        RECT 54.000 103.600 54.800 104.400 ;
        RECT 54.100 100.400 54.700 103.600 ;
        RECT 54.000 99.600 54.800 100.400 ;
        RECT 55.700 98.400 56.300 105.600 ;
        RECT 54.000 97.600 54.800 98.400 ;
        RECT 55.600 97.600 56.400 98.400 ;
        RECT 46.000 93.600 46.800 94.400 ;
        RECT 47.600 93.600 48.400 94.400 ;
        RECT 46.100 92.400 46.700 93.600 ;
        RECT 44.400 91.600 45.200 92.400 ;
        RECT 46.000 91.600 46.800 92.400 ;
        RECT 38.000 87.600 38.800 88.400 ;
        RECT 28.400 83.600 29.200 84.400 ;
        RECT 44.500 82.400 45.100 91.600 ;
        RECT 46.000 88.300 46.800 88.400 ;
        RECT 47.700 88.300 48.300 93.600 ;
        RECT 46.000 87.700 48.300 88.300 ;
        RECT 54.100 88.300 54.700 97.600 ;
        RECT 55.600 91.600 56.400 92.400 ;
        RECT 55.700 90.400 56.300 91.600 ;
        RECT 55.600 89.600 56.400 90.400 ;
        RECT 57.300 88.400 57.900 107.600 ;
        RECT 66.900 102.400 67.500 107.600 ;
        RECT 71.700 106.400 72.300 107.600 ;
        RECT 78.100 106.400 78.700 107.600 ;
        RECT 71.600 105.600 72.400 106.400 ;
        RECT 78.000 105.600 78.800 106.400 ;
        RECT 79.600 105.600 80.400 106.400 ;
        RECT 73.200 103.600 74.000 104.400 ;
        RECT 63.600 101.600 64.400 102.400 ;
        RECT 66.800 101.600 67.600 102.400 ;
        RECT 71.600 101.600 72.400 102.400 ;
        RECT 60.400 93.600 61.200 94.400 ;
        RECT 58.800 89.600 59.600 90.400 ;
        RECT 55.600 88.300 56.400 88.400 ;
        RECT 54.100 87.700 56.400 88.300 ;
        RECT 46.000 87.600 46.800 87.700 ;
        RECT 55.600 87.600 56.400 87.700 ;
        RECT 57.200 87.600 58.000 88.400 ;
        RECT 57.200 83.600 58.000 84.400 ;
        RECT 44.400 81.600 45.200 82.400 ;
        RECT 44.500 78.400 45.100 81.600 ;
        RECT 57.300 80.400 57.900 83.600 ;
        RECT 57.200 79.600 58.000 80.400 ;
        RECT 44.400 77.600 45.200 78.400 ;
        RECT 31.600 75.600 32.400 76.400 ;
        RECT 30.000 73.600 30.800 74.400 ;
        RECT 26.800 67.600 27.600 68.400 ;
        RECT 23.600 61.600 24.400 62.400 ;
        RECT 20.500 59.700 22.700 60.300 ;
        RECT 20.500 58.400 21.100 59.700 ;
        RECT 30.100 58.400 30.700 73.600 ;
        RECT 31.700 72.400 32.300 75.600 ;
        RECT 58.900 74.400 59.500 89.600 ;
        RECT 60.500 78.400 61.100 93.600 ;
        RECT 63.700 90.400 64.300 101.600 ;
        RECT 71.700 98.400 72.300 101.600 ;
        RECT 71.600 97.600 72.400 98.400 ;
        RECT 68.400 95.600 69.200 96.400 ;
        RECT 66.800 91.600 67.600 92.400 ;
        RECT 62.000 89.600 62.800 90.400 ;
        RECT 63.600 89.600 64.400 90.400 ;
        RECT 68.500 88.400 69.100 95.600 ;
        RECT 73.300 92.400 73.900 103.600 ;
        RECT 73.200 91.600 74.000 92.400 ;
        RECT 78.000 91.600 78.800 92.400 ;
        RECT 68.400 87.600 69.200 88.400 ;
        RECT 78.100 86.400 78.700 91.600 ;
        RECT 78.000 85.600 78.800 86.400 ;
        RECT 66.800 83.600 67.600 84.400 ;
        RECT 62.000 79.600 62.800 80.400 ;
        RECT 60.400 77.600 61.200 78.400 ;
        RECT 60.400 75.600 61.200 76.400 ;
        RECT 58.800 73.600 59.600 74.400 ;
        RECT 31.600 71.600 32.400 72.400 ;
        RECT 33.200 71.600 34.000 72.400 ;
        RECT 36.400 71.800 37.200 72.600 ;
        RECT 43.000 71.800 43.800 72.600 ;
        RECT 31.600 69.600 32.400 70.400 ;
        RECT 31.700 62.400 32.300 69.600 ;
        RECT 31.600 61.600 32.400 62.400 ;
        RECT 12.400 57.600 13.200 58.400 ;
        RECT 20.400 57.600 21.200 58.400 ;
        RECT 30.000 57.600 30.800 58.400 ;
        RECT 33.300 56.400 33.900 71.600 ;
        RECT 36.400 68.400 37.000 71.800 ;
        RECT 40.400 68.400 41.200 68.600 ;
        RECT 36.400 67.800 41.200 68.400 ;
        RECT 36.400 67.000 37.000 67.800 ;
        RECT 37.800 67.000 38.600 67.200 ;
        RECT 41.200 67.000 42.000 67.200 ;
        RECT 43.200 67.000 43.800 71.800 ;
        RECT 46.000 71.600 46.800 72.400 ;
        RECT 54.000 71.600 54.800 72.400 ;
        RECT 36.400 66.200 37.200 67.000 ;
        RECT 37.800 66.400 42.000 67.000 ;
        RECT 43.000 66.200 43.800 67.000 ;
        RECT 41.200 63.600 42.000 64.400 ;
        RECT 41.200 61.600 42.000 62.400 ;
        RECT 15.600 55.600 16.400 56.400 ;
        RECT 15.700 54.400 16.300 55.600 ;
        RECT 23.600 55.000 24.400 55.800 ;
        RECT 25.000 55.000 29.200 55.600 ;
        RECT 30.200 55.000 31.000 55.800 ;
        RECT 33.200 55.600 34.000 56.400 ;
        RECT 38.000 55.600 38.800 56.400 ;
        RECT 15.600 53.600 16.400 54.400 ;
        RECT 23.600 54.200 24.200 55.000 ;
        RECT 25.000 54.800 25.800 55.000 ;
        RECT 28.400 54.800 29.200 55.000 ;
        RECT 23.600 53.600 28.400 54.200 ;
        RECT 10.800 51.600 11.600 52.400 ;
        RECT 17.200 51.600 18.000 52.400 ;
        RECT 10.900 50.400 11.500 51.600 ;
        RECT 10.800 49.600 11.600 50.400 ;
        RECT 23.600 50.200 24.200 53.600 ;
        RECT 27.600 53.400 28.400 53.600 ;
        RECT 30.400 50.200 31.000 55.000 ;
        RECT 31.600 53.600 32.400 54.400 ;
        RECT 31.700 52.400 32.300 53.600 ;
        RECT 31.600 51.600 32.400 52.400 ;
        RECT 23.600 49.400 24.400 50.200 ;
        RECT 30.200 49.400 31.000 50.200 ;
        RECT 22.000 47.600 22.800 48.400 ;
        RECT 22.100 38.400 22.700 47.600 ;
        RECT 25.200 43.600 26.000 44.400 ;
        RECT 22.000 37.600 22.800 38.400 ;
        RECT 25.300 32.400 25.900 43.600 ;
        RECT 38.100 38.400 38.700 55.600 ;
        RECT 41.300 54.400 41.900 61.600 ;
        RECT 42.800 57.600 43.600 58.400 ;
        RECT 41.200 53.600 42.000 54.400 ;
        RECT 42.900 52.400 43.500 57.600 ;
        RECT 39.600 51.600 40.400 52.400 ;
        RECT 42.800 51.600 43.600 52.400 ;
        RECT 41.200 45.600 42.000 46.400 ;
        RECT 38.000 37.600 38.800 38.400 ;
        RECT 41.300 36.400 41.900 45.600 ;
        RECT 31.600 35.600 32.400 36.400 ;
        RECT 41.200 35.600 42.000 36.400 ;
        RECT 31.700 34.400 32.300 35.600 ;
        RECT 31.600 33.600 32.400 34.400 ;
        RECT 34.800 33.600 35.600 34.400 ;
        RECT 34.900 32.400 35.500 33.600 ;
        RECT 9.200 31.600 10.000 32.400 ;
        RECT 25.200 31.600 26.000 32.400 ;
        RECT 34.800 31.600 35.600 32.400 ;
        RECT 7.600 29.600 8.400 30.400 ;
        RECT 9.300 28.400 9.900 31.600 ;
        RECT 41.300 30.400 41.900 35.600 ;
        RECT 46.100 34.400 46.700 71.600 ;
        RECT 54.100 70.400 54.700 71.600 ;
        RECT 54.000 69.600 54.800 70.400 ;
        RECT 58.800 69.600 59.600 70.400 ;
        RECT 60.500 68.400 61.100 75.600 ;
        RECT 62.100 70.400 62.700 79.600 ;
        RECT 63.600 77.600 64.400 78.400 ;
        RECT 63.700 70.400 64.300 77.600 ;
        RECT 66.900 76.400 67.500 83.600 ;
        RECT 66.800 75.600 67.600 76.400 ;
        RECT 66.800 73.600 67.600 74.400 ;
        RECT 70.000 73.600 70.800 74.400 ;
        RECT 66.900 72.400 67.500 73.600 ;
        RECT 70.100 72.400 70.700 73.600 ;
        RECT 79.700 72.400 80.300 105.600 ;
        RECT 66.800 71.600 67.600 72.400 ;
        RECT 70.000 71.600 70.800 72.400 ;
        RECT 73.200 72.300 74.000 72.400 ;
        RECT 71.700 71.700 74.000 72.300 ;
        RECT 62.000 69.600 62.800 70.400 ;
        RECT 63.600 69.600 64.400 70.400 ;
        RECT 65.200 69.600 66.000 70.400 ;
        RECT 68.400 69.600 69.200 70.400 ;
        RECT 71.700 68.400 72.300 71.700 ;
        RECT 73.200 71.600 74.000 71.700 ;
        RECT 79.600 71.600 80.400 72.400 ;
        RECT 60.400 67.600 61.200 68.400 ;
        RECT 68.400 67.600 69.200 68.400 ;
        RECT 71.600 67.600 72.400 68.400 ;
        RECT 73.200 67.600 74.000 68.400 ;
        RECT 76.400 67.600 77.200 68.400 ;
        RECT 79.600 67.600 80.400 68.400 ;
        RECT 81.300 68.300 81.900 123.600 ;
        RECT 86.100 114.400 86.700 131.600 ;
        RECT 86.000 113.600 86.800 114.400 ;
        RECT 86.100 108.400 86.700 113.600 ;
        RECT 84.400 107.600 85.200 108.400 ;
        RECT 86.000 107.600 86.800 108.400 ;
        RECT 86.000 96.300 86.800 96.400 ;
        RECT 87.700 96.300 88.300 133.600 ;
        RECT 95.700 118.400 96.300 133.600 ;
        RECT 97.000 130.200 97.600 135.000 ;
        RECT 98.800 134.800 99.600 135.000 ;
        RECT 102.200 134.800 103.000 135.000 ;
        RECT 103.800 134.200 104.400 135.000 ;
        RECT 99.600 133.600 104.400 134.200 ;
        RECT 119.600 133.600 120.400 134.400 ;
        RECT 122.800 133.600 123.600 134.400 ;
        RECT 99.600 133.400 100.400 133.600 ;
        RECT 102.000 131.600 102.800 132.400 ;
        RECT 103.800 130.200 104.400 133.600 ;
        RECT 119.700 132.400 120.300 133.600 ;
        RECT 110.000 131.600 110.800 132.400 ;
        RECT 119.600 131.600 120.400 132.400 ;
        RECT 121.200 131.600 122.000 132.400 ;
        RECT 97.000 129.400 97.800 130.200 ;
        RECT 103.600 129.400 104.400 130.200 ;
        RECT 95.600 117.600 96.400 118.400 ;
        RECT 101.800 111.800 102.600 112.600 ;
        RECT 108.400 111.800 109.200 112.600 ;
        RECT 95.600 109.600 96.400 110.400 ;
        RECT 92.400 107.600 93.200 108.400 ;
        RECT 95.600 107.600 96.400 108.400 ;
        RECT 100.400 107.600 101.200 108.400 ;
        RECT 90.800 105.600 91.600 106.400 ;
        RECT 92.500 98.400 93.100 107.600 ;
        RECT 95.700 98.400 96.300 107.600 ;
        RECT 100.500 104.300 101.100 107.600 ;
        RECT 101.800 107.000 102.400 111.800 ;
        RECT 104.400 108.400 105.200 108.600 ;
        RECT 108.600 108.400 109.200 111.800 ;
        RECT 104.400 107.800 109.200 108.400 ;
        RECT 103.600 107.000 104.400 107.200 ;
        RECT 107.000 107.000 107.800 107.200 ;
        RECT 108.600 107.000 109.200 107.800 ;
        RECT 101.800 106.200 102.600 107.000 ;
        RECT 103.600 106.400 107.800 107.000 ;
        RECT 108.400 106.200 109.200 107.000 ;
        RECT 100.500 103.700 102.700 104.300 ;
        RECT 102.100 98.400 102.700 103.700 ;
        RECT 92.400 97.600 93.200 98.400 ;
        RECT 95.600 97.600 96.400 98.400 ;
        RECT 102.000 97.600 102.800 98.400 ;
        RECT 86.000 95.700 88.300 96.300 ;
        RECT 86.000 95.600 86.800 95.700 ;
        RECT 86.000 93.600 86.800 94.400 ;
        RECT 90.800 93.600 91.600 94.400 ;
        RECT 90.900 92.400 91.500 93.600 ;
        RECT 87.600 91.600 88.400 92.400 ;
        RECT 90.800 91.600 91.600 92.400 ;
        RECT 86.000 83.600 86.800 84.400 ;
        RECT 82.800 75.600 83.600 76.400 ;
        RECT 84.400 73.600 85.200 74.400 ;
        RECT 84.500 70.400 85.100 73.600 ;
        RECT 86.100 72.400 86.700 83.600 ;
        RECT 87.600 77.600 88.400 78.400 ;
        RECT 86.000 71.600 86.800 72.400 ;
        RECT 87.700 70.400 88.300 77.600 ;
        RECT 89.200 75.600 90.000 76.400 ;
        RECT 89.300 74.400 89.900 75.600 ;
        RECT 89.200 73.600 90.000 74.400 ;
        RECT 84.400 69.600 85.200 70.400 ;
        RECT 87.600 69.600 88.400 70.400 ;
        RECT 90.900 68.400 91.500 91.600 ;
        RECT 92.500 78.400 93.100 97.600 ;
        RECT 95.600 95.600 96.400 96.400 ;
        RECT 95.700 80.400 96.300 95.600 ;
        RECT 108.400 93.600 109.200 94.400 ;
        RECT 108.500 92.400 109.100 93.600 ;
        RECT 97.200 91.600 98.000 92.400 ;
        RECT 108.400 91.600 109.200 92.400 ;
        RECT 97.300 90.400 97.900 91.600 ;
        RECT 97.200 89.600 98.000 90.400 ;
        RECT 105.200 89.600 106.000 90.400 ;
        RECT 110.100 82.400 110.700 131.600 ;
        RECT 113.200 129.600 114.000 130.400 ;
        RECT 111.600 123.600 112.400 124.400 ;
        RECT 111.700 110.400 112.300 123.600 ;
        RECT 113.300 118.400 113.900 129.600 ;
        RECT 113.200 117.600 114.000 118.400 ;
        RECT 121.300 110.400 121.900 131.600 ;
        RECT 111.600 109.600 112.400 110.400 ;
        RECT 113.200 109.600 114.000 110.400 ;
        RECT 121.200 109.600 122.000 110.400 ;
        RECT 111.700 108.400 112.300 109.600 ;
        RECT 113.300 108.400 113.900 109.600 ;
        RECT 111.600 107.600 112.400 108.400 ;
        RECT 113.200 107.600 114.000 108.400 ;
        RECT 119.600 107.600 120.400 108.400 ;
        RECT 118.000 105.600 118.800 106.400 ;
        RECT 121.300 106.300 121.900 109.600 ;
        RECT 124.500 106.400 125.100 135.600 ;
        RECT 127.600 131.600 128.400 132.400 ;
        RECT 130.800 131.600 131.600 132.400 ;
        RECT 137.200 131.600 138.000 132.400 ;
        RECT 146.800 131.600 147.600 132.400 ;
        RECT 130.900 118.400 131.500 131.600 ;
        RECT 137.300 130.400 137.900 131.600 ;
        RECT 137.200 129.600 138.000 130.400 ;
        RECT 175.600 123.600 176.400 124.400 ;
        RECT 130.800 117.600 131.600 118.400 ;
        RECT 145.200 111.400 146.000 112.400 ;
        RECT 154.800 111.600 155.600 112.400 ;
        RECT 166.000 111.600 166.800 112.400 ;
        RECT 154.900 110.400 155.500 111.600 ;
        RECT 166.100 110.400 166.700 111.600 ;
        RECT 175.700 110.400 176.300 123.600 ;
        RECT 135.600 109.600 136.400 110.400 ;
        RECT 148.400 109.600 149.200 110.400 ;
        RECT 154.800 109.600 155.600 110.400 ;
        RECT 162.800 109.600 163.600 110.400 ;
        RECT 166.000 109.600 166.800 110.400 ;
        RECT 175.600 109.600 176.400 110.400 ;
        RECT 137.200 107.600 138.000 108.400 ;
        RECT 150.000 107.600 150.800 108.400 ;
        RECT 158.000 107.600 158.800 108.400 ;
        RECT 164.400 107.600 165.200 108.400 ;
        RECT 170.800 107.600 171.600 108.400 ;
        RECT 119.700 105.700 121.900 106.300 ;
        RECT 118.100 100.400 118.700 105.600 ;
        RECT 118.000 99.600 118.800 100.400 ;
        RECT 119.700 98.400 120.300 105.700 ;
        RECT 124.400 105.600 125.200 106.400 ;
        RECT 135.600 105.600 136.400 106.400 ;
        RECT 137.300 98.400 137.900 107.600 ;
        RECT 150.100 106.400 150.700 107.600 ;
        RECT 148.400 105.600 149.200 106.400 ;
        RECT 150.000 105.600 150.800 106.400 ;
        RECT 166.000 105.600 166.800 106.400 ;
        RECT 154.800 103.600 155.600 104.400 ;
        RECT 159.600 103.600 160.400 104.400 ;
        RECT 119.600 97.600 120.400 98.400 ;
        RECT 137.200 97.600 138.000 98.400 ;
        RECT 111.600 95.600 112.400 96.400 ;
        RECT 132.600 95.600 133.400 95.800 ;
        RECT 111.700 94.400 112.300 95.600 ;
        RECT 132.600 95.000 138.200 95.600 ;
        RECT 138.800 95.000 139.600 95.800 ;
        RECT 143.600 95.600 144.400 96.400 ;
        RECT 111.600 93.600 112.400 94.400 ;
        RECT 114.800 93.600 115.600 94.400 ;
        RECT 121.200 93.600 122.000 94.400 ;
        RECT 111.700 92.400 112.300 93.600 ;
        RECT 114.900 92.400 115.500 93.600 ;
        RECT 111.600 91.600 112.400 92.400 ;
        RECT 114.800 91.600 115.600 92.400 ;
        RECT 116.400 91.600 117.200 92.400 ;
        RECT 113.200 89.600 114.000 90.400 ;
        RECT 110.000 81.600 110.800 82.400 ;
        RECT 95.600 79.600 96.400 80.400 ;
        RECT 110.000 79.600 110.800 80.400 ;
        RECT 92.400 77.600 93.200 78.400 ;
        RECT 106.800 73.600 107.600 74.400 ;
        RECT 94.000 71.600 94.800 72.400 ;
        RECT 97.200 71.800 98.000 72.600 ;
        RECT 103.400 71.800 104.200 72.600 ;
        RECT 106.900 72.400 107.500 73.600 ;
        RECT 82.800 68.300 83.600 68.400 ;
        RECT 81.300 67.700 83.600 68.300 ;
        RECT 82.800 67.600 83.600 67.700 ;
        RECT 84.400 67.600 85.200 68.400 ;
        RECT 90.800 67.600 91.600 68.400 ;
        RECT 57.200 65.600 58.000 66.400 ;
        RECT 57.300 64.400 57.900 65.600 ;
        RECT 57.200 63.600 58.000 64.400 ;
        RECT 68.500 58.400 69.100 67.600 ;
        RECT 73.200 63.600 74.000 64.400 ;
        RECT 68.400 57.600 69.200 58.400 ;
        RECT 73.300 56.400 73.900 63.600 ;
        RECT 76.400 57.600 77.200 58.400 ;
        RECT 76.500 56.400 77.100 57.600 ;
        RECT 73.200 55.600 74.000 56.400 ;
        RECT 76.400 55.600 77.200 56.400 ;
        RECT 54.000 53.600 54.800 54.400 ;
        RECT 54.100 52.400 54.700 53.600 ;
        RECT 54.000 51.600 54.800 52.400 ;
        RECT 55.600 51.600 56.400 52.400 ;
        RECT 65.200 51.600 66.000 52.400 ;
        RECT 73.200 51.600 74.000 52.400 ;
        RECT 74.800 51.600 75.600 52.400 ;
        RECT 55.700 48.400 56.300 51.600 ;
        RECT 65.300 50.400 65.900 51.600 ;
        RECT 63.600 49.600 64.400 50.400 ;
        RECT 65.200 49.600 66.000 50.400 ;
        RECT 68.400 49.600 69.200 50.400 ;
        RECT 55.600 47.600 56.400 48.400 ;
        RECT 54.000 45.600 54.800 46.400 ;
        RECT 63.700 44.400 64.300 49.600 ;
        RECT 66.800 45.600 67.600 46.400 ;
        RECT 63.600 43.600 64.400 44.400 ;
        RECT 65.200 41.600 66.000 42.400 ;
        RECT 46.000 33.600 46.800 34.400 ;
        RECT 42.800 31.600 43.600 32.400 ;
        RECT 44.200 31.800 45.000 32.600 ;
        RECT 50.800 31.800 51.600 32.600 ;
        RECT 15.600 29.600 16.400 30.400 ;
        RECT 22.000 29.600 22.800 30.400 ;
        RECT 39.600 29.600 40.400 30.400 ;
        RECT 41.200 29.600 42.000 30.400 ;
        RECT 9.200 27.600 10.000 28.400 ;
        RECT 10.800 25.600 11.600 26.400 ;
        RECT 4.400 23.600 5.200 24.400 ;
        RECT 4.500 12.400 5.100 23.600 ;
        RECT 10.900 18.400 11.500 25.600 ;
        RECT 14.000 23.600 14.800 24.400 ;
        RECT 10.800 17.600 11.600 18.400 ;
        RECT 14.100 14.400 14.700 23.600 ;
        RECT 15.700 14.400 16.300 29.600 ;
        RECT 22.100 28.400 22.700 29.600 ;
        RECT 39.700 28.400 40.300 29.600 ;
        RECT 42.900 28.400 43.500 31.600 ;
        RECT 17.200 27.600 18.000 28.400 ;
        RECT 20.400 27.600 21.200 28.400 ;
        RECT 22.000 27.600 22.800 28.400 ;
        RECT 38.000 27.600 38.800 28.400 ;
        RECT 39.600 27.600 40.400 28.400 ;
        RECT 42.800 27.600 43.600 28.400 ;
        RECT 20.500 26.400 21.100 27.600 ;
        RECT 44.200 27.000 44.800 31.800 ;
        RECT 46.800 28.400 47.600 28.600 ;
        RECT 51.000 28.400 51.600 31.800 ;
        RECT 65.300 30.400 65.900 41.600 ;
        RECT 65.200 29.600 66.000 30.400 ;
        RECT 46.800 27.800 51.600 28.400 ;
        RECT 46.000 27.000 46.800 27.200 ;
        RECT 49.400 27.000 50.200 27.200 ;
        RECT 51.000 27.000 51.600 27.800 ;
        RECT 20.400 25.600 21.200 26.400 ;
        RECT 26.800 25.600 27.600 26.400 ;
        RECT 44.200 26.200 45.000 27.000 ;
        RECT 46.000 26.400 50.200 27.000 ;
        RECT 50.800 26.200 51.600 27.000 ;
        RECT 46.000 23.600 46.800 24.400 ;
        RECT 57.200 23.600 58.000 24.400 ;
        RECT 25.200 17.600 26.000 18.400 ;
        RECT 26.800 17.600 27.600 18.400 ;
        RECT 42.800 17.600 43.600 18.400 ;
        RECT 44.400 17.600 45.200 18.400 ;
        RECT 14.000 13.600 14.800 14.400 ;
        RECT 15.600 13.600 16.400 14.400 ;
        RECT 22.000 13.600 22.800 14.400 ;
        RECT 15.700 12.400 16.300 13.600 ;
        RECT 25.300 12.400 25.900 17.600 ;
        RECT 26.900 16.400 27.500 17.600 ;
        RECT 26.800 15.600 27.600 16.400 ;
        RECT 42.900 16.300 43.500 17.600 ;
        RECT 44.500 16.400 45.100 17.600 ;
        RECT 41.300 15.700 43.500 16.300 ;
        RECT 41.300 12.400 41.900 15.700 ;
        RECT 44.400 15.600 45.200 16.400 ;
        RECT 46.100 14.400 46.700 23.600 ;
        RECT 42.800 13.600 43.600 14.400 ;
        RECT 46.000 13.600 46.800 14.400 ;
        RECT 57.300 12.400 57.900 23.600 ;
        RECT 66.900 18.400 67.500 45.600 ;
        RECT 70.000 43.600 70.800 44.400 ;
        RECT 70.100 28.400 70.700 43.600 ;
        RECT 70.000 27.600 70.800 28.400 ;
        RECT 68.400 25.600 69.200 26.400 ;
        RECT 68.500 18.400 69.100 25.600 ;
        RECT 73.300 18.400 73.900 51.600 ;
        RECT 79.700 48.400 80.300 67.600 ;
        RECT 81.200 63.600 82.000 64.400 ;
        RECT 81.300 52.400 81.900 63.600 ;
        RECT 84.500 58.400 85.100 67.600 ;
        RECT 94.100 66.400 94.700 71.600 ;
        RECT 97.200 68.400 97.800 71.800 ;
        RECT 102.200 69.800 103.000 70.600 ;
        RECT 102.200 68.400 102.800 69.800 ;
        RECT 97.200 67.800 102.800 68.400 ;
        RECT 97.200 67.000 97.800 67.800 ;
        RECT 98.600 67.000 99.400 67.200 ;
        RECT 102.000 67.000 102.800 67.200 ;
        RECT 103.600 67.000 104.200 71.800 ;
        RECT 106.800 71.600 107.600 72.400 ;
        RECT 110.100 70.400 110.700 79.600 ;
        RECT 113.300 78.400 113.900 89.600 ;
        RECT 114.800 83.600 115.600 84.400 ;
        RECT 113.200 77.600 114.000 78.400 ;
        RECT 110.000 69.600 110.800 70.400 ;
        RECT 111.600 67.600 112.400 68.400 ;
        RECT 94.000 65.600 94.800 66.400 ;
        RECT 97.200 66.200 98.000 67.000 ;
        RECT 98.600 66.400 104.200 67.000 ;
        RECT 103.400 66.200 104.200 66.400 ;
        RECT 89.200 63.600 90.000 64.400 ;
        RECT 92.400 63.600 93.200 64.400 ;
        RECT 98.800 63.600 99.600 64.400 ;
        RECT 84.400 57.600 85.200 58.400 ;
        RECT 86.000 53.600 86.800 54.400 ;
        RECT 86.100 52.400 86.700 53.600 ;
        RECT 81.200 51.600 82.000 52.400 ;
        RECT 86.000 51.600 86.800 52.400 ;
        RECT 82.800 49.600 83.600 50.400 ;
        RECT 79.600 47.600 80.400 48.400 ;
        RECT 82.900 46.400 83.500 49.600 ;
        RECT 82.800 45.600 83.600 46.400 ;
        RECT 78.000 43.600 78.800 44.400 ;
        RECT 74.800 35.600 75.600 36.400 ;
        RECT 74.900 28.400 75.500 35.600 ;
        RECT 76.400 31.600 77.200 32.400 ;
        RECT 76.400 29.600 77.200 30.400 ;
        RECT 76.500 28.400 77.100 29.600 ;
        RECT 74.800 27.600 75.600 28.400 ;
        RECT 76.400 27.600 77.200 28.400 ;
        RECT 66.800 17.600 67.600 18.400 ;
        RECT 68.400 17.600 69.200 18.400 ;
        RECT 73.200 17.600 74.000 18.400 ;
        RECT 71.600 15.600 72.400 16.400 ;
        RECT 76.400 15.600 77.200 16.400 ;
        RECT 71.700 14.400 72.300 15.600 ;
        RECT 76.500 14.400 77.100 15.600 ;
        RECT 78.100 14.400 78.700 43.600 ;
        RECT 92.500 36.400 93.100 63.600 ;
        RECT 97.200 59.600 98.000 60.400 ;
        RECT 95.600 57.600 96.400 58.400 ;
        RECT 92.400 35.600 93.200 36.400 ;
        RECT 79.600 31.600 80.400 32.400 ;
        RECT 82.800 31.800 83.600 32.600 ;
        RECT 89.400 31.800 90.200 32.600 ;
        RECT 79.700 30.400 80.300 31.600 ;
        RECT 79.600 29.600 80.400 30.400 ;
        RECT 82.800 28.400 83.400 31.800 ;
        RECT 86.800 28.400 87.600 28.600 ;
        RECT 81.200 27.600 82.000 28.400 ;
        RECT 82.800 27.800 87.600 28.400 ;
        RECT 82.800 27.000 83.400 27.800 ;
        RECT 84.200 27.000 85.000 27.200 ;
        RECT 87.600 27.000 88.400 27.200 ;
        RECT 89.600 27.000 90.200 31.800 ;
        RECT 95.700 30.400 96.300 57.600 ;
        RECT 97.300 56.400 97.900 59.600 ;
        RECT 97.200 55.600 98.000 56.400 ;
        RECT 98.900 54.400 99.500 63.600 ;
        RECT 111.700 58.400 112.300 67.600 ;
        RECT 113.200 63.600 114.000 64.400 ;
        RECT 113.300 58.400 113.900 63.600 ;
        RECT 111.600 57.600 112.400 58.400 ;
        RECT 113.200 57.600 114.000 58.400 ;
        RECT 110.000 55.600 110.800 56.400 ;
        RECT 113.200 55.600 114.000 56.400 ;
        RECT 114.900 56.300 115.500 83.600 ;
        RECT 116.500 64.400 117.100 91.600 ;
        RECT 121.300 90.400 121.900 93.600 ;
        RECT 124.400 91.600 125.200 92.400 ;
        RECT 124.500 90.400 125.100 91.600 ;
        RECT 121.200 89.600 122.000 90.400 ;
        RECT 124.400 89.600 125.200 90.400 ;
        RECT 132.600 90.200 133.200 95.000 ;
        RECT 134.000 94.800 134.800 95.000 ;
        RECT 137.400 94.800 138.200 95.000 ;
        RECT 139.000 94.200 139.600 95.000 ;
        RECT 143.700 94.400 144.300 95.600 ;
        RECT 134.000 93.600 139.600 94.200 ;
        RECT 143.600 93.600 144.400 94.400 ;
        RECT 148.400 93.600 149.200 94.400 ;
        RECT 153.200 93.600 154.000 94.400 ;
        RECT 134.000 92.200 134.600 93.600 ;
        RECT 133.800 91.400 134.600 92.200 ;
        RECT 139.000 90.200 139.600 93.600 ;
        RECT 145.200 91.600 146.000 92.400 ;
        RECT 132.600 89.400 133.400 90.200 ;
        RECT 138.800 89.400 139.600 90.200 ;
        RECT 142.000 89.600 142.800 90.400 ;
        RECT 148.400 89.600 149.200 90.400 ;
        RECT 142.100 84.400 142.700 89.600 ;
        RECT 153.300 84.400 153.900 93.600 ;
        RECT 154.900 92.400 155.500 103.600 ;
        RECT 158.000 94.300 158.800 94.400 ;
        RECT 159.700 94.300 160.300 103.600 ;
        RECT 166.100 98.400 166.700 105.600 ;
        RECT 166.000 97.600 166.800 98.400 ;
        RECT 162.800 95.600 163.600 96.400 ;
        RECT 164.600 95.600 165.400 95.800 ;
        RECT 162.900 94.400 163.500 95.600 ;
        RECT 164.600 95.000 170.200 95.600 ;
        RECT 170.800 95.000 171.600 95.800 ;
        RECT 158.000 93.700 160.300 94.300 ;
        RECT 158.000 93.600 158.800 93.700 ;
        RECT 162.800 93.600 163.600 94.400 ;
        RECT 154.800 91.600 155.600 92.400 ;
        RECT 158.100 90.400 158.700 93.600 ;
        RECT 158.000 89.600 158.800 90.400 ;
        RECT 161.200 89.600 162.000 90.400 ;
        RECT 162.800 89.600 163.600 90.400 ;
        RECT 164.600 90.200 165.200 95.000 ;
        RECT 166.000 94.800 166.800 95.000 ;
        RECT 169.400 94.800 170.200 95.000 ;
        RECT 171.000 94.200 171.600 95.000 ;
        RECT 166.000 93.600 171.600 94.200 ;
        RECT 166.000 92.200 166.600 93.600 ;
        RECT 165.800 91.400 166.600 92.200 ;
        RECT 171.000 90.200 171.600 93.600 ;
        RECT 121.200 83.600 122.000 84.400 ;
        RECT 142.000 83.600 142.800 84.400 ;
        RECT 153.200 83.600 154.000 84.400 ;
        RECT 154.800 83.600 155.600 84.400 ;
        RECT 159.600 83.600 160.400 84.400 ;
        RECT 119.600 81.600 120.400 82.400 ;
        RECT 116.400 63.600 117.200 64.400 ;
        RECT 116.500 58.400 117.100 63.600 ;
        RECT 116.400 57.600 117.200 58.400 ;
        RECT 119.700 56.400 120.300 81.600 ;
        RECT 121.300 78.400 121.900 83.600 ;
        RECT 121.200 77.600 122.000 78.400 ;
        RECT 130.800 73.600 131.600 74.400 ;
        RECT 142.000 73.600 142.800 74.400 ;
        RECT 142.100 72.400 142.700 73.600 ;
        RECT 140.400 71.600 141.200 72.400 ;
        RECT 142.000 71.600 142.800 72.400 ;
        RECT 145.200 71.600 146.000 72.400 ;
        RECT 150.200 71.800 151.000 72.600 ;
        RECT 154.900 72.400 155.500 83.600 ;
        RECT 159.700 80.400 160.300 83.600 ;
        RECT 159.600 79.600 160.400 80.400 ;
        RECT 145.300 70.400 145.900 71.600 ;
        RECT 145.200 69.600 146.000 70.400 ;
        RECT 132.400 67.600 133.200 68.400 ;
        RECT 137.200 68.300 138.000 68.400 ;
        RECT 137.200 67.700 139.500 68.300 ;
        RECT 137.200 67.600 138.000 67.700 ;
        RECT 132.500 66.400 133.100 67.600 ;
        RECT 132.400 65.600 133.200 66.400 ;
        RECT 121.200 63.600 122.000 64.400 ;
        RECT 114.900 55.700 117.100 56.300 ;
        RECT 110.100 54.400 110.700 55.600 ;
        RECT 98.800 53.600 99.600 54.400 ;
        RECT 100.400 53.600 101.200 54.400 ;
        RECT 110.000 53.600 110.800 54.400 ;
        RECT 113.300 54.300 113.900 55.600 ;
        RECT 116.500 54.400 117.100 55.700 ;
        RECT 119.600 55.600 120.400 56.400 ;
        RECT 119.700 54.400 120.300 55.600 ;
        RECT 114.800 54.300 115.600 54.400 ;
        RECT 113.300 53.700 115.600 54.300 ;
        RECT 114.800 53.600 115.600 53.700 ;
        RECT 116.400 53.600 117.200 54.400 ;
        RECT 119.600 53.600 120.400 54.400 ;
        RECT 97.200 51.600 98.000 52.400 ;
        RECT 97.300 48.400 97.900 51.600 ;
        RECT 100.500 50.400 101.100 53.600 ;
        RECT 103.600 51.600 104.400 52.400 ;
        RECT 108.400 51.600 109.200 52.400 ;
        RECT 111.600 51.600 112.400 52.400 ;
        RECT 111.700 50.400 112.300 51.600 ;
        RECT 116.500 50.400 117.100 53.600 ;
        RECT 121.300 50.400 121.900 63.600 ;
        RECT 124.400 57.600 125.200 58.400 ;
        RECT 124.500 52.400 125.100 57.600 ;
        RECT 124.400 51.600 125.200 52.400 ;
        RECT 100.400 49.600 101.200 50.400 ;
        RECT 111.600 49.600 112.400 50.400 ;
        RECT 113.200 49.600 114.000 50.400 ;
        RECT 116.400 49.600 117.200 50.400 ;
        RECT 121.200 49.600 122.000 50.400 ;
        RECT 97.200 47.600 98.000 48.400 ;
        RECT 97.300 42.400 97.900 47.600 ;
        RECT 102.000 43.600 102.800 44.400 ;
        RECT 97.200 41.600 98.000 42.400 ;
        RECT 102.100 32.400 102.700 43.600 ;
        RECT 111.700 38.400 112.300 49.600 ;
        RECT 111.600 37.600 112.400 38.400 ;
        RECT 105.200 33.600 106.000 34.400 ;
        RECT 105.300 32.400 105.900 33.600 ;
        RECT 102.000 31.600 102.800 32.400 ;
        RECT 105.200 31.600 106.000 32.400 ;
        RECT 106.800 31.600 107.600 32.400 ;
        RECT 111.600 31.600 112.400 32.400 ;
        RECT 102.100 30.400 102.700 31.600 ;
        RECT 105.300 30.400 105.900 31.600 ;
        RECT 106.900 30.400 107.500 31.600 ;
        RECT 113.300 30.400 113.900 49.600 ;
        RECT 121.200 47.600 122.000 48.400 ;
        RECT 118.000 43.600 118.800 44.400 ;
        RECT 116.400 32.300 117.200 32.400 ;
        RECT 118.100 32.300 118.700 43.600 ;
        RECT 119.600 37.600 120.400 38.400 ;
        RECT 132.500 32.400 133.100 65.600 ;
        RECT 138.900 56.400 139.500 67.700 ;
        RECT 143.600 67.600 144.400 68.400 ;
        RECT 148.400 67.600 149.200 68.400 ;
        RECT 150.200 67.000 150.800 71.800 ;
        RECT 154.800 71.600 155.600 72.400 ;
        RECT 156.400 71.800 157.200 72.600 ;
        RECT 151.400 69.800 152.200 70.600 ;
        RECT 151.600 68.400 152.200 69.800 ;
        RECT 156.600 68.400 157.200 71.800 ;
        RECT 151.600 67.800 157.200 68.400 ;
        RECT 151.600 67.000 152.400 67.200 ;
        RECT 155.000 67.000 155.800 67.200 ;
        RECT 156.600 67.000 157.200 67.800 ;
        RECT 161.300 68.300 161.900 89.600 ;
        RECT 162.900 78.400 163.500 89.600 ;
        RECT 164.600 89.400 165.400 90.200 ;
        RECT 170.800 89.400 171.600 90.200 ;
        RECT 175.600 83.600 176.400 84.400 ;
        RECT 162.800 77.600 163.600 78.400 ;
        RECT 161.300 67.700 163.500 68.300 ;
        RECT 150.200 66.400 155.800 67.000 ;
        RECT 150.200 66.200 151.000 66.400 ;
        RECT 156.400 66.200 157.200 67.000 ;
        RECT 140.400 63.600 141.200 64.400 ;
        RECT 154.800 63.600 155.600 64.400 ;
        RECT 161.200 63.600 162.000 64.400 ;
        RECT 138.800 55.600 139.600 56.400 ;
        RECT 140.500 54.400 141.100 63.600 ;
        RECT 142.200 55.600 143.000 55.800 ;
        RECT 142.200 55.000 147.800 55.600 ;
        RECT 148.400 55.000 149.200 55.800 ;
        RECT 134.000 53.600 134.800 54.400 ;
        RECT 138.800 53.600 139.600 54.400 ;
        RECT 140.400 53.600 141.200 54.400 ;
        RECT 134.100 52.400 134.700 53.600 ;
        RECT 134.000 51.600 134.800 52.400 ;
        RECT 135.600 51.600 136.400 52.400 ;
        RECT 140.400 51.600 141.200 52.400 ;
        RECT 135.700 48.400 136.300 51.600 ;
        RECT 134.000 47.600 134.800 48.400 ;
        RECT 135.600 47.600 136.400 48.400 ;
        RECT 116.400 31.700 118.700 32.300 ;
        RECT 116.400 31.600 117.200 31.700 ;
        RECT 118.100 30.400 118.700 31.700 ;
        RECT 132.400 31.600 133.200 32.400 ;
        RECT 90.800 29.600 91.600 30.400 ;
        RECT 95.600 29.600 96.400 30.400 ;
        RECT 102.000 29.600 102.800 30.400 ;
        RECT 103.600 29.600 104.400 30.400 ;
        RECT 105.200 29.600 106.000 30.400 ;
        RECT 106.800 29.600 107.600 30.400 ;
        RECT 113.200 29.600 114.000 30.400 ;
        RECT 118.000 29.600 118.800 30.400 ;
        RECT 129.200 29.600 130.000 30.400 ;
        RECT 90.900 28.400 91.500 29.600 ;
        RECT 113.300 28.400 113.900 29.600 ;
        RECT 90.800 27.600 91.600 28.400 ;
        RECT 110.000 27.600 110.800 28.400 ;
        RECT 113.200 27.600 114.000 28.400 ;
        RECT 82.800 26.200 83.600 27.000 ;
        RECT 84.200 26.400 88.400 27.000 ;
        RECT 89.400 26.200 90.200 27.000 ;
        RECT 97.200 25.600 98.000 26.400 ;
        RECT 87.600 23.600 88.400 24.400 ;
        RECT 86.000 17.600 86.800 18.400 ;
        RECT 71.600 13.600 72.400 14.400 ;
        RECT 76.400 13.600 77.200 14.400 ;
        RECT 78.000 13.600 78.800 14.400 ;
        RECT 86.100 12.400 86.700 17.600 ;
        RECT 87.700 14.400 88.300 23.600 ;
        RECT 97.300 18.400 97.900 25.600 ;
        RECT 89.200 17.600 90.000 18.400 ;
        RECT 97.200 17.600 98.000 18.400 ;
        RECT 106.800 17.600 107.600 18.400 ;
        RECT 89.300 16.400 89.900 17.600 ;
        RECT 97.300 16.400 97.900 17.600 ;
        RECT 89.200 15.600 90.000 16.400 ;
        RECT 97.200 15.600 98.000 16.400 ;
        RECT 102.000 15.000 102.800 15.800 ;
        RECT 108.200 15.600 109.000 15.800 ;
        RECT 103.400 15.000 109.000 15.600 ;
        RECT 87.600 13.600 88.400 14.400 ;
        RECT 102.000 14.200 102.600 15.000 ;
        RECT 103.400 14.800 104.200 15.000 ;
        RECT 106.800 14.800 107.600 15.000 ;
        RECT 102.000 13.600 107.600 14.200 ;
        RECT 4.400 11.600 5.200 12.400 ;
        RECT 14.000 11.600 14.800 12.400 ;
        RECT 15.600 11.600 16.400 12.400 ;
        RECT 25.200 11.600 26.000 12.400 ;
        RECT 26.800 11.600 27.600 12.400 ;
        RECT 41.200 11.600 42.000 12.400 ;
        RECT 44.400 11.600 45.200 12.400 ;
        RECT 57.200 11.600 58.000 12.400 ;
        RECT 63.600 11.600 64.400 12.400 ;
        RECT 70.000 11.600 70.800 12.400 ;
        RECT 73.200 11.600 74.000 12.400 ;
        RECT 84.400 11.600 85.200 12.400 ;
        RECT 86.000 11.600 86.800 12.400 ;
        RECT 73.300 10.400 73.900 11.600 ;
        RECT 73.200 9.600 74.000 10.400 ;
        RECT 102.000 10.200 102.600 13.600 ;
        RECT 107.000 12.200 107.600 13.600 ;
        RECT 107.000 11.400 107.800 12.200 ;
        RECT 108.400 10.200 109.000 15.000 ;
        RECT 110.100 14.400 110.700 27.600 ;
        RECT 114.800 23.600 115.600 24.400 ;
        RECT 114.900 18.400 115.500 23.600 ;
        RECT 111.600 17.600 112.400 18.400 ;
        RECT 114.800 17.600 115.600 18.400 ;
        RECT 111.700 14.400 112.300 17.600 ;
        RECT 113.400 15.600 114.200 15.800 ;
        RECT 113.400 15.000 119.000 15.600 ;
        RECT 119.600 15.000 120.400 15.800 ;
        RECT 110.000 13.600 110.800 14.400 ;
        RECT 111.600 13.600 112.400 14.400 ;
        RECT 102.000 9.400 102.800 10.200 ;
        RECT 108.200 9.400 109.000 10.200 ;
        RECT 113.400 10.200 114.000 15.000 ;
        RECT 114.800 14.800 115.600 15.000 ;
        RECT 118.200 14.800 119.000 15.000 ;
        RECT 119.800 14.200 120.400 15.000 ;
        RECT 114.800 13.600 120.400 14.200 ;
        RECT 129.200 13.600 130.000 14.400 ;
        RECT 132.400 13.600 133.200 14.400 ;
        RECT 114.800 12.200 115.400 13.600 ;
        RECT 114.600 11.400 115.400 12.200 ;
        RECT 119.800 10.200 120.400 13.600 ;
        RECT 129.300 12.400 129.900 13.600 ;
        RECT 132.500 12.400 133.100 13.600 ;
        RECT 134.100 12.400 134.700 47.600 ;
        RECT 140.500 30.400 141.100 51.600 ;
        RECT 142.200 50.200 142.800 55.000 ;
        RECT 143.600 54.800 144.400 55.000 ;
        RECT 147.000 54.800 147.800 55.000 ;
        RECT 148.600 54.200 149.200 55.000 ;
        RECT 154.900 54.400 155.500 63.600 ;
        RECT 156.400 56.300 157.200 56.400 ;
        RECT 156.400 55.700 158.700 56.300 ;
        RECT 156.400 55.600 157.200 55.700 ;
        RECT 143.600 53.600 149.200 54.200 ;
        RECT 154.800 53.600 155.600 54.400 ;
        RECT 143.600 52.200 144.200 53.600 ;
        RECT 143.400 51.400 144.200 52.200 ;
        RECT 148.600 50.200 149.200 53.600 ;
        RECT 156.400 51.600 157.200 52.400 ;
        RECT 142.200 49.400 143.000 50.200 ;
        RECT 148.400 49.400 149.200 50.200 ;
        RECT 143.600 43.600 144.400 44.400 ;
        RECT 140.400 29.600 141.200 30.400 ;
        RECT 143.700 28.400 144.300 43.600 ;
        RECT 148.600 31.800 149.400 32.600 ;
        RECT 154.800 31.800 155.600 32.600 ;
        RECT 135.600 27.600 136.400 28.400 ;
        RECT 143.600 27.600 144.400 28.400 ;
        RECT 146.800 27.600 147.600 28.400 ;
        RECT 148.600 27.000 149.200 31.800 ;
        RECT 149.800 29.800 150.600 30.600 ;
        RECT 150.000 28.400 150.600 29.800 ;
        RECT 155.000 28.400 155.600 31.800 ;
        RECT 150.000 27.800 155.600 28.400 ;
        RECT 150.000 27.000 150.800 27.200 ;
        RECT 153.400 27.000 154.200 27.200 ;
        RECT 155.000 27.000 155.600 27.800 ;
        RECT 148.600 26.400 154.200 27.000 ;
        RECT 140.400 25.600 141.200 26.400 ;
        RECT 148.600 26.200 149.400 26.400 ;
        RECT 154.800 26.200 155.600 27.000 ;
        RECT 140.500 24.400 141.100 25.600 ;
        RECT 158.100 24.400 158.700 55.700 ;
        RECT 161.300 52.400 161.900 63.600 ;
        RECT 161.200 51.600 162.000 52.400 ;
        RECT 161.200 49.600 162.000 50.400 ;
        RECT 162.900 46.400 163.500 67.700 ;
        RECT 175.700 58.400 176.300 83.600 ;
        RECT 175.600 57.600 176.400 58.400 ;
        RECT 164.400 53.600 165.200 54.400 ;
        RECT 164.500 52.400 165.100 53.600 ;
        RECT 164.400 51.600 165.200 52.400 ;
        RECT 169.200 51.600 170.000 52.400 ;
        RECT 169.300 50.400 169.900 51.600 ;
        RECT 169.200 49.600 170.000 50.400 ;
        RECT 162.800 45.600 163.600 46.400 ;
        RECT 167.600 45.600 168.400 46.400 ;
        RECT 161.200 29.600 162.000 30.400 ;
        RECT 162.800 29.600 163.600 30.400 ;
        RECT 159.600 25.600 160.400 26.400 ;
        RECT 159.700 24.400 160.300 25.600 ;
        RECT 135.600 23.600 136.400 24.400 ;
        RECT 140.400 23.600 141.200 24.400 ;
        RECT 142.000 23.600 142.800 24.400 ;
        RECT 158.000 23.600 158.800 24.400 ;
        RECT 159.600 23.600 160.400 24.400 ;
        RECT 135.700 16.400 136.300 23.600 ;
        RECT 135.600 15.600 136.400 16.400 ;
        RECT 135.600 13.600 136.400 14.400 ;
        RECT 142.100 12.400 142.700 23.600 ;
        RECT 158.100 16.400 158.700 23.600 ;
        RECT 158.000 15.600 158.800 16.400 ;
        RECT 159.600 15.600 160.400 16.400 ;
        RECT 159.700 14.400 160.300 15.600 ;
        RECT 154.800 13.600 155.600 14.400 ;
        RECT 159.600 13.600 160.400 14.400 ;
        RECT 154.900 12.400 155.500 13.600 ;
        RECT 161.300 12.400 161.900 29.600 ;
        RECT 167.700 18.400 168.300 45.600 ;
        RECT 175.600 43.600 176.400 44.400 ;
        RECT 169.200 23.600 170.000 24.400 ;
        RECT 170.800 23.600 171.600 24.400 ;
        RECT 169.300 22.400 169.900 23.600 ;
        RECT 169.200 21.600 170.000 22.400 ;
        RECT 167.600 17.600 168.400 18.400 ;
        RECT 170.900 12.400 171.500 23.600 ;
        RECT 175.700 14.400 176.300 43.600 ;
        RECT 177.200 21.600 178.000 22.400 ;
        RECT 172.400 13.600 173.200 14.400 ;
        RECT 175.600 13.600 176.400 14.400 ;
        RECT 177.300 12.400 177.900 21.600 ;
        RECT 129.200 11.600 130.000 12.400 ;
        RECT 132.400 11.600 133.200 12.400 ;
        RECT 134.000 11.600 134.800 12.400 ;
        RECT 140.400 11.600 141.200 12.400 ;
        RECT 142.000 11.600 142.800 12.400 ;
        RECT 145.200 11.600 146.000 12.400 ;
        RECT 154.800 11.600 155.600 12.400 ;
        RECT 161.200 11.600 162.000 12.400 ;
        RECT 162.800 11.600 163.600 12.400 ;
        RECT 170.800 11.600 171.600 12.400 ;
        RECT 177.200 11.600 178.000 12.400 ;
        RECT 113.400 9.400 114.200 10.200 ;
        RECT 119.600 9.400 120.400 10.200 ;
      LAYER via2 ;
        RECT 145.200 111.600 146.000 112.400 ;
      LAYER metal3 ;
        RECT 74.800 138.300 75.600 138.400 ;
        RECT 30.100 137.700 75.600 138.300 ;
        RECT 30.100 136.400 30.700 137.700 ;
        RECT 74.800 137.600 75.600 137.700 ;
        RECT 20.400 136.300 21.200 136.400 ;
        RECT 30.000 136.300 30.800 136.400 ;
        RECT 20.400 135.700 30.800 136.300 ;
        RECT 20.400 135.600 21.200 135.700 ;
        RECT 30.000 135.600 30.800 135.700 ;
        RECT 49.200 136.300 50.000 136.400 ;
        RECT 62.000 136.300 62.800 136.400 ;
        RECT 49.200 135.700 62.800 136.300 ;
        RECT 49.200 135.600 50.000 135.700 ;
        RECT 62.000 135.600 62.800 135.700 ;
        RECT 78.000 134.300 78.800 134.400 ;
        RECT 74.900 133.700 78.800 134.300 ;
        RECT 9.200 132.300 10.000 132.400 ;
        RECT 12.400 132.300 13.200 132.400 ;
        RECT 9.200 131.700 13.200 132.300 ;
        RECT 9.200 131.600 10.000 131.700 ;
        RECT 12.400 131.600 13.200 131.700 ;
        RECT 17.200 132.300 18.000 132.400 ;
        RECT 28.400 132.300 29.200 132.400 ;
        RECT 17.200 131.700 29.200 132.300 ;
        RECT 17.200 131.600 18.000 131.700 ;
        RECT 28.400 131.600 29.200 131.700 ;
        RECT 33.200 132.300 34.000 132.400 ;
        RECT 49.200 132.300 50.000 132.400 ;
        RECT 33.200 131.700 50.000 132.300 ;
        RECT 33.200 131.600 34.000 131.700 ;
        RECT 49.200 131.600 50.000 131.700 ;
        RECT 60.400 132.300 61.200 132.400 ;
        RECT 74.900 132.300 75.500 133.700 ;
        RECT 78.000 133.600 78.800 133.700 ;
        RECT 82.800 134.300 83.600 134.400 ;
        RECT 90.800 134.300 91.600 134.400 ;
        RECT 122.800 134.300 123.600 134.400 ;
        RECT 82.800 133.700 91.600 134.300 ;
        RECT 82.800 133.600 83.600 133.700 ;
        RECT 90.800 133.600 91.600 133.700 ;
        RECT 118.100 133.700 123.600 134.300 ;
        RECT 60.400 131.700 75.500 132.300 ;
        RECT 76.400 132.300 77.200 132.400 ;
        RECT 86.000 132.300 86.800 132.400 ;
        RECT 76.400 131.700 86.800 132.300 ;
        RECT 60.400 131.600 61.200 131.700 ;
        RECT 76.400 131.600 77.200 131.700 ;
        RECT 86.000 131.600 86.800 131.700 ;
        RECT 102.000 132.300 102.800 132.400 ;
        RECT 118.100 132.300 118.700 133.700 ;
        RECT 122.800 133.600 123.600 133.700 ;
        RECT 102.000 131.700 118.700 132.300 ;
        RECT 119.600 132.300 120.400 132.400 ;
        RECT 127.600 132.300 128.400 132.400 ;
        RECT 119.600 131.700 128.400 132.300 ;
        RECT 102.000 131.600 102.800 131.700 ;
        RECT 119.600 131.600 120.400 131.700 ;
        RECT 127.600 131.600 128.400 131.700 ;
        RECT 130.800 132.300 131.600 132.400 ;
        RECT 146.800 132.300 147.600 132.400 ;
        RECT 130.800 131.700 147.600 132.300 ;
        RECT 130.800 131.600 131.600 131.700 ;
        RECT 146.800 131.600 147.600 131.700 ;
        RECT 23.600 130.300 24.400 130.400 ;
        RECT 34.800 130.300 35.600 130.400 ;
        RECT 23.600 129.700 35.600 130.300 ;
        RECT 23.600 129.600 24.400 129.700 ;
        RECT 34.800 129.600 35.600 129.700 ;
        RECT 73.200 130.300 74.000 130.400 ;
        RECT 79.600 130.300 80.400 130.400 ;
        RECT 73.200 129.700 80.400 130.300 ;
        RECT 73.200 129.600 74.000 129.700 ;
        RECT 79.600 129.600 80.400 129.700 ;
        RECT 113.200 130.300 114.000 130.400 ;
        RECT 137.200 130.300 138.000 130.400 ;
        RECT 113.200 129.700 138.000 130.300 ;
        RECT 113.200 129.600 114.000 129.700 ;
        RECT 137.200 129.600 138.000 129.700 ;
        RECT 10.800 128.300 11.600 128.400 ;
        RECT 23.700 128.300 24.300 129.600 ;
        RECT 10.800 127.700 24.300 128.300 ;
        RECT 28.400 128.300 29.200 128.400 ;
        RECT 38.000 128.300 38.800 128.400 ;
        RECT 62.000 128.300 62.800 128.400 ;
        RECT 28.400 127.700 62.800 128.300 ;
        RECT 10.800 127.600 11.600 127.700 ;
        RECT 28.400 127.600 29.200 127.700 ;
        RECT 38.000 127.600 38.800 127.700 ;
        RECT 62.000 127.600 62.800 127.700 ;
        RECT 68.400 128.300 69.200 128.400 ;
        RECT 84.400 128.300 85.200 128.400 ;
        RECT 68.400 127.700 85.200 128.300 ;
        RECT 68.400 127.600 69.200 127.700 ;
        RECT 84.400 127.600 85.200 127.700 ;
        RECT 34.800 114.300 35.600 114.400 ;
        RECT 42.800 114.300 43.600 114.400 ;
        RECT 34.800 113.700 43.600 114.300 ;
        RECT 34.800 113.600 35.600 113.700 ;
        RECT 42.800 113.600 43.600 113.700 ;
        RECT 60.400 114.300 61.200 114.400 ;
        RECT 86.000 114.300 86.800 114.400 ;
        RECT 60.400 113.700 86.800 114.300 ;
        RECT 60.400 113.600 61.200 113.700 ;
        RECT 86.000 113.600 86.800 113.700 ;
        RECT 6.000 112.300 6.800 112.400 ;
        RECT 22.000 112.300 22.800 112.400 ;
        RECT 6.000 111.700 22.800 112.300 ;
        RECT 6.000 111.600 6.800 111.700 ;
        RECT 22.000 111.600 22.800 111.700 ;
        RECT 62.000 112.300 62.800 112.400 ;
        RECT 70.000 112.300 70.800 112.400 ;
        RECT 62.000 111.700 70.800 112.300 ;
        RECT 62.000 111.600 62.800 111.700 ;
        RECT 70.000 111.600 70.800 111.700 ;
        RECT 145.200 112.300 146.000 112.400 ;
        RECT 166.000 112.300 166.800 112.400 ;
        RECT 145.200 111.700 166.800 112.300 ;
        RECT 145.200 111.600 146.000 111.700 ;
        RECT 166.000 111.600 166.800 111.700 ;
        RECT 52.400 110.300 53.200 110.400 ;
        RECT 60.400 110.300 61.200 110.400 ;
        RECT 52.400 109.700 61.200 110.300 ;
        RECT 52.400 109.600 53.200 109.700 ;
        RECT 60.400 109.600 61.200 109.700 ;
        RECT 76.400 110.300 77.200 110.400 ;
        RECT 79.600 110.300 80.400 110.400 ;
        RECT 76.400 109.700 80.400 110.300 ;
        RECT 76.400 109.600 77.200 109.700 ;
        RECT 79.600 109.600 80.400 109.700 ;
        RECT 95.600 110.300 96.400 110.400 ;
        RECT 111.600 110.300 112.400 110.400 ;
        RECT 95.600 109.700 112.400 110.300 ;
        RECT 95.600 109.600 96.400 109.700 ;
        RECT 111.600 109.600 112.400 109.700 ;
        RECT 121.200 110.300 122.000 110.400 ;
        RECT 135.600 110.300 136.400 110.400 ;
        RECT 148.400 110.300 149.200 110.400 ;
        RECT 121.200 109.700 149.200 110.300 ;
        RECT 121.200 109.600 122.000 109.700 ;
        RECT 135.600 109.600 136.400 109.700 ;
        RECT 148.400 109.600 149.200 109.700 ;
        RECT 154.800 110.300 155.600 110.400 ;
        RECT 162.800 110.300 163.600 110.400 ;
        RECT 175.600 110.300 176.400 110.400 ;
        RECT 154.800 109.700 176.400 110.300 ;
        RECT 154.800 109.600 155.600 109.700 ;
        RECT 162.800 109.600 163.600 109.700 ;
        RECT 175.600 109.600 176.400 109.700 ;
        RECT 12.400 108.300 13.200 108.400 ;
        RECT 18.800 108.300 19.600 108.400 ;
        RECT 12.400 107.700 19.600 108.300 ;
        RECT 12.400 107.600 13.200 107.700 ;
        RECT 18.800 107.600 19.600 107.700 ;
        RECT 44.400 108.300 45.200 108.400 ;
        RECT 58.800 108.300 59.600 108.400 ;
        RECT 44.400 107.700 59.600 108.300 ;
        RECT 44.400 107.600 45.200 107.700 ;
        RECT 58.800 107.600 59.600 107.700 ;
        RECT 65.200 108.300 66.000 108.400 ;
        RECT 84.400 108.300 85.200 108.400 ;
        RECT 65.200 107.700 85.200 108.300 ;
        RECT 65.200 107.600 66.000 107.700 ;
        RECT 84.400 107.600 85.200 107.700 ;
        RECT 86.000 108.300 86.800 108.400 ;
        RECT 95.600 108.300 96.400 108.400 ;
        RECT 86.000 107.700 96.400 108.300 ;
        RECT 86.000 107.600 86.800 107.700 ;
        RECT 95.600 107.600 96.400 107.700 ;
        RECT 113.200 108.300 114.000 108.400 ;
        RECT 119.600 108.300 120.400 108.400 ;
        RECT 113.200 107.700 120.400 108.300 ;
        RECT 113.200 107.600 114.000 107.700 ;
        RECT 119.600 107.600 120.400 107.700 ;
        RECT 158.000 108.300 158.800 108.400 ;
        RECT 164.400 108.300 165.200 108.400 ;
        RECT 170.800 108.300 171.600 108.400 ;
        RECT 158.000 107.700 171.600 108.300 ;
        RECT 158.000 107.600 158.800 107.700 ;
        RECT 164.400 107.600 165.200 107.700 ;
        RECT 170.800 107.600 171.600 107.700 ;
        RECT 2.800 106.300 3.600 106.400 ;
        RECT 10.800 106.300 11.600 106.400 ;
        RECT 2.800 105.700 11.600 106.300 ;
        RECT 2.800 105.600 3.600 105.700 ;
        RECT 10.800 105.600 11.600 105.700 ;
        RECT 15.600 106.300 16.400 106.400 ;
        RECT 39.600 106.300 40.400 106.400 ;
        RECT 15.600 105.700 40.400 106.300 ;
        RECT 15.600 105.600 16.400 105.700 ;
        RECT 39.600 105.600 40.400 105.700 ;
        RECT 42.800 106.300 43.600 106.400 ;
        RECT 50.800 106.300 51.600 106.400 ;
        RECT 42.800 105.700 51.600 106.300 ;
        RECT 42.800 105.600 43.600 105.700 ;
        RECT 50.800 105.600 51.600 105.700 ;
        RECT 71.600 106.300 72.400 106.400 ;
        RECT 78.000 106.300 78.800 106.400 ;
        RECT 90.800 106.300 91.600 106.400 ;
        RECT 71.600 105.700 91.600 106.300 ;
        RECT 71.600 105.600 72.400 105.700 ;
        RECT 78.000 105.600 78.800 105.700 ;
        RECT 90.800 105.600 91.600 105.700 ;
        RECT 124.400 106.300 125.200 106.400 ;
        RECT 135.600 106.300 136.400 106.400 ;
        RECT 148.400 106.300 149.200 106.400 ;
        RECT 124.400 105.700 149.200 106.300 ;
        RECT 124.400 105.600 125.200 105.700 ;
        RECT 135.600 105.600 136.400 105.700 ;
        RECT 148.400 105.600 149.200 105.700 ;
        RECT 150.000 106.300 150.800 106.400 ;
        RECT 166.000 106.300 166.800 106.400 ;
        RECT 150.000 105.700 166.800 106.300 ;
        RECT 150.000 105.600 150.800 105.700 ;
        RECT 166.000 105.600 166.800 105.700 ;
        RECT 10.900 104.300 11.500 105.600 ;
        RECT 18.800 104.300 19.600 104.400 ;
        RECT 20.400 104.300 21.200 104.400 ;
        RECT 10.900 103.700 21.200 104.300 ;
        RECT 18.800 103.600 19.600 103.700 ;
        RECT 20.400 103.600 21.200 103.700 ;
        RECT 25.200 102.300 26.000 102.400 ;
        RECT 63.600 102.300 64.400 102.400 ;
        RECT 25.200 101.700 64.400 102.300 ;
        RECT 25.200 101.600 26.000 101.700 ;
        RECT 63.600 101.600 64.400 101.700 ;
        RECT 66.800 102.300 67.600 102.400 ;
        RECT 71.600 102.300 72.400 102.400 ;
        RECT 66.800 101.700 72.400 102.300 ;
        RECT 66.800 101.600 67.600 101.700 ;
        RECT 71.600 101.600 72.400 101.700 ;
        RECT 54.000 100.300 54.800 100.400 ;
        RECT 97.200 100.300 98.000 100.400 ;
        RECT 118.000 100.300 118.800 100.400 ;
        RECT 54.000 99.700 118.800 100.300 ;
        RECT 54.000 99.600 54.800 99.700 ;
        RECT 97.200 99.600 98.000 99.700 ;
        RECT 118.000 99.600 118.800 99.700 ;
        RECT 33.200 98.300 34.000 98.400 ;
        RECT 54.000 98.300 54.800 98.400 ;
        RECT 33.200 97.700 54.800 98.300 ;
        RECT 33.200 97.600 34.000 97.700 ;
        RECT 54.000 97.600 54.800 97.700 ;
        RECT 55.600 98.300 56.400 98.400 ;
        RECT 92.400 98.300 93.200 98.400 ;
        RECT 55.600 97.700 93.200 98.300 ;
        RECT 55.600 97.600 56.400 97.700 ;
        RECT 92.400 97.600 93.200 97.700 ;
        RECT 4.400 95.600 5.200 96.400 ;
        RECT 68.400 96.300 69.200 96.400 ;
        RECT 86.000 96.300 86.800 96.400 ;
        RECT 68.400 95.700 86.800 96.300 ;
        RECT 68.400 95.600 69.200 95.700 ;
        RECT 86.000 95.600 86.800 95.700 ;
        RECT 143.600 96.300 144.400 96.400 ;
        RECT 162.800 96.300 163.600 96.400 ;
        RECT 143.600 95.700 163.600 96.300 ;
        RECT 143.600 95.600 144.400 95.700 ;
        RECT 162.800 95.600 163.600 95.700 ;
        RECT 7.600 94.300 8.400 94.400 ;
        RECT 22.000 94.300 22.800 94.400 ;
        RECT 7.600 93.700 22.800 94.300 ;
        RECT 7.600 93.600 8.400 93.700 ;
        RECT 22.000 93.600 22.800 93.700 ;
        RECT 25.200 94.300 26.000 94.400 ;
        RECT 28.400 94.300 29.200 94.400 ;
        RECT 25.200 93.700 29.200 94.300 ;
        RECT 25.200 93.600 26.000 93.700 ;
        RECT 28.400 93.600 29.200 93.700 ;
        RECT 47.600 94.300 48.400 94.400 ;
        RECT 86.000 94.300 86.800 94.400 ;
        RECT 47.600 93.700 86.800 94.300 ;
        RECT 47.600 93.600 48.400 93.700 ;
        RECT 86.000 93.600 86.800 93.700 ;
        RECT 108.400 94.300 109.200 94.400 ;
        RECT 114.800 94.300 115.600 94.400 ;
        RECT 148.400 94.300 149.200 94.400 ;
        RECT 108.400 93.700 149.200 94.300 ;
        RECT 108.400 93.600 109.200 93.700 ;
        RECT 114.800 93.600 115.600 93.700 ;
        RECT 148.400 93.600 149.200 93.700 ;
        RECT 17.200 92.300 18.000 92.400 ;
        RECT 20.400 92.300 21.200 92.400 ;
        RECT 46.000 92.300 46.800 92.400 ;
        RECT 17.200 91.700 46.800 92.300 ;
        RECT 17.200 91.600 18.000 91.700 ;
        RECT 20.400 91.600 21.200 91.700 ;
        RECT 46.000 91.600 46.800 91.700 ;
        RECT 66.800 92.300 67.600 92.400 ;
        RECT 73.200 92.300 74.000 92.400 ;
        RECT 66.800 91.700 74.000 92.300 ;
        RECT 66.800 91.600 67.600 91.700 ;
        RECT 73.200 91.600 74.000 91.700 ;
        RECT 87.600 92.300 88.400 92.400 ;
        RECT 90.800 92.300 91.600 92.400 ;
        RECT 87.600 91.700 91.600 92.300 ;
        RECT 87.600 91.600 88.400 91.700 ;
        RECT 90.800 91.600 91.600 91.700 ;
        RECT 111.600 92.300 112.400 92.400 ;
        RECT 124.400 92.300 125.200 92.400 ;
        RECT 145.200 92.300 146.000 92.400 ;
        RECT 154.800 92.300 155.600 92.400 ;
        RECT 111.600 91.700 155.600 92.300 ;
        RECT 111.600 91.600 112.400 91.700 ;
        RECT 124.400 91.600 125.200 91.700 ;
        RECT 145.200 91.600 146.000 91.700 ;
        RECT 154.800 91.600 155.600 91.700 ;
        RECT 15.600 90.300 16.400 90.400 ;
        RECT 23.600 90.300 24.400 90.400 ;
        RECT 15.600 89.700 24.400 90.300 ;
        RECT 15.600 89.600 16.400 89.700 ;
        RECT 23.600 89.600 24.400 89.700 ;
        RECT 34.800 90.300 35.600 90.400 ;
        RECT 55.600 90.300 56.400 90.400 ;
        RECT 34.800 89.700 56.400 90.300 ;
        RECT 34.800 89.600 35.600 89.700 ;
        RECT 55.600 89.600 56.400 89.700 ;
        RECT 62.000 90.300 62.800 90.400 ;
        RECT 97.200 90.300 98.000 90.400 ;
        RECT 62.000 89.700 98.000 90.300 ;
        RECT 62.000 89.600 62.800 89.700 ;
        RECT 97.200 89.600 98.000 89.700 ;
        RECT 105.200 90.300 106.000 90.400 ;
        RECT 113.200 90.300 114.000 90.400 ;
        RECT 121.200 90.300 122.000 90.400 ;
        RECT 105.200 89.700 122.000 90.300 ;
        RECT 105.200 89.600 106.000 89.700 ;
        RECT 113.200 89.600 114.000 89.700 ;
        RECT 121.200 89.600 122.000 89.700 ;
        RECT 148.400 90.300 149.200 90.400 ;
        RECT 162.800 90.300 163.600 90.400 ;
        RECT 148.400 89.700 163.600 90.300 ;
        RECT 148.400 89.600 149.200 89.700 ;
        RECT 162.800 89.600 163.600 89.700 ;
        RECT 18.800 88.300 19.600 88.400 ;
        RECT 38.000 88.300 38.800 88.400 ;
        RECT 18.800 87.700 38.800 88.300 ;
        RECT 18.800 87.600 19.600 87.700 ;
        RECT 38.000 87.600 38.800 87.700 ;
        RECT 57.200 88.300 58.000 88.400 ;
        RECT 68.400 88.300 69.200 88.400 ;
        RECT 57.200 87.700 69.200 88.300 ;
        RECT 57.200 87.600 58.000 87.700 ;
        RECT 68.400 87.600 69.200 87.700 ;
        RECT 38.100 86.300 38.700 87.600 ;
        RECT 78.000 86.300 78.800 86.400 ;
        RECT 38.100 85.700 78.800 86.300 ;
        RECT 78.000 85.600 78.800 85.700 ;
        RECT 28.400 84.300 29.200 84.400 ;
        RECT 86.000 84.300 86.800 84.400 ;
        RECT 28.400 83.700 86.800 84.300 ;
        RECT 28.400 83.600 29.200 83.700 ;
        RECT 86.000 83.600 86.800 83.700 ;
        RECT 121.200 84.300 122.000 84.400 ;
        RECT 142.000 84.300 142.800 84.400 ;
        RECT 121.200 83.700 142.800 84.300 ;
        RECT 121.200 83.600 122.000 83.700 ;
        RECT 142.000 83.600 142.800 83.700 ;
        RECT 153.200 84.300 154.000 84.400 ;
        RECT 175.600 84.300 176.400 84.400 ;
        RECT 153.200 83.700 176.400 84.300 ;
        RECT 153.200 83.600 154.000 83.700 ;
        RECT 175.600 83.600 176.400 83.700 ;
        RECT 22.000 82.300 22.800 82.400 ;
        RECT 44.400 82.300 45.200 82.400 ;
        RECT 22.000 81.700 45.200 82.300 ;
        RECT 22.000 81.600 22.800 81.700 ;
        RECT 44.400 81.600 45.200 81.700 ;
        RECT 110.000 82.300 110.800 82.400 ;
        RECT 119.600 82.300 120.400 82.400 ;
        RECT 110.000 81.700 120.400 82.300 ;
        RECT 110.000 81.600 110.800 81.700 ;
        RECT 119.600 81.600 120.400 81.700 ;
        RECT 57.200 80.300 58.000 80.400 ;
        RECT 62.000 80.300 62.800 80.400 ;
        RECT 57.200 79.700 62.800 80.300 ;
        RECT 57.200 79.600 58.000 79.700 ;
        RECT 62.000 79.600 62.800 79.700 ;
        RECT 95.600 80.300 96.400 80.400 ;
        RECT 110.000 80.300 110.800 80.400 ;
        RECT 159.600 80.300 160.400 80.400 ;
        RECT 95.600 79.700 160.400 80.300 ;
        RECT 95.600 79.600 96.400 79.700 ;
        RECT 110.000 79.600 110.800 79.700 ;
        RECT 159.600 79.600 160.400 79.700 ;
        RECT 44.400 78.300 45.200 78.400 ;
        RECT 60.400 78.300 61.200 78.400 ;
        RECT 44.400 77.700 61.200 78.300 ;
        RECT 44.400 77.600 45.200 77.700 ;
        RECT 60.400 77.600 61.200 77.700 ;
        RECT 63.600 78.300 64.400 78.400 ;
        RECT 87.600 78.300 88.400 78.400 ;
        RECT 63.600 77.700 88.400 78.300 ;
        RECT 63.600 77.600 64.400 77.700 ;
        RECT 87.600 77.600 88.400 77.700 ;
        RECT 60.400 76.300 61.200 76.400 ;
        RECT 66.800 76.300 67.600 76.400 ;
        RECT 60.400 75.700 67.600 76.300 ;
        RECT 60.400 75.600 61.200 75.700 ;
        RECT 66.800 75.600 67.600 75.700 ;
        RECT 82.800 76.300 83.600 76.400 ;
        RECT 89.200 76.300 90.000 76.400 ;
        RECT 82.800 75.700 90.000 76.300 ;
        RECT 82.800 75.600 83.600 75.700 ;
        RECT 89.200 75.600 90.000 75.700 ;
        RECT 7.600 74.300 8.400 74.400 ;
        RECT 17.200 74.300 18.000 74.400 ;
        RECT 7.600 73.700 18.000 74.300 ;
        RECT 7.600 73.600 8.400 73.700 ;
        RECT 17.200 73.600 18.000 73.700 ;
        RECT 18.800 74.300 19.600 74.400 ;
        RECT 25.200 74.300 26.000 74.400 ;
        RECT 30.000 74.300 30.800 74.400 ;
        RECT 18.800 73.700 30.800 74.300 ;
        RECT 18.800 73.600 19.600 73.700 ;
        RECT 25.200 73.600 26.000 73.700 ;
        RECT 30.000 73.600 30.800 73.700 ;
        RECT 58.800 74.300 59.600 74.400 ;
        RECT 66.800 74.300 67.600 74.400 ;
        RECT 84.400 74.300 85.200 74.400 ;
        RECT 106.800 74.300 107.600 74.400 ;
        RECT 130.800 74.300 131.600 74.400 ;
        RECT 142.000 74.300 142.800 74.400 ;
        RECT 58.800 73.700 142.800 74.300 ;
        RECT 58.800 73.600 59.600 73.700 ;
        RECT 66.800 73.600 67.600 73.700 ;
        RECT 84.400 73.600 85.200 73.700 ;
        RECT 106.800 73.600 107.600 73.700 ;
        RECT 130.800 73.600 131.600 73.700 ;
        RECT 142.000 73.600 142.800 73.700 ;
        RECT 4.400 72.300 5.200 72.400 ;
        RECT 6.000 72.300 6.800 72.400 ;
        RECT 4.400 71.700 6.800 72.300 ;
        RECT 4.400 71.600 5.200 71.700 ;
        RECT 6.000 71.600 6.800 71.700 ;
        RECT 31.600 72.300 32.400 72.400 ;
        RECT 54.000 72.300 54.800 72.400 ;
        RECT 70.000 72.300 70.800 72.400 ;
        RECT 31.600 71.700 70.800 72.300 ;
        RECT 31.600 71.600 32.400 71.700 ;
        RECT 54.000 71.600 54.800 71.700 ;
        RECT 70.000 71.600 70.800 71.700 ;
        RECT 78.000 72.300 78.800 72.400 ;
        RECT 79.600 72.300 80.400 72.400 ;
        RECT 94.000 72.300 94.800 72.400 ;
        RECT 78.000 71.700 94.800 72.300 ;
        RECT 78.000 71.600 78.800 71.700 ;
        RECT 79.600 71.600 80.400 71.700 ;
        RECT 94.000 71.600 94.800 71.700 ;
        RECT 140.400 72.300 141.200 72.400 ;
        RECT 145.200 72.300 146.000 72.400 ;
        RECT 154.800 72.300 155.600 72.400 ;
        RECT 140.400 71.700 155.600 72.300 ;
        RECT 140.400 71.600 141.200 71.700 ;
        RECT 145.200 71.600 146.000 71.700 ;
        RECT 154.800 71.600 155.600 71.700 ;
        RECT 58.800 70.300 59.600 70.400 ;
        RECT 63.600 70.300 64.400 70.400 ;
        RECT 58.800 69.700 64.400 70.300 ;
        RECT 58.800 69.600 59.600 69.700 ;
        RECT 63.600 69.600 64.400 69.700 ;
        RECT 65.200 70.300 66.000 70.400 ;
        RECT 68.400 70.300 69.200 70.400 ;
        RECT 65.200 69.700 69.200 70.300 ;
        RECT 65.200 69.600 66.000 69.700 ;
        RECT 68.400 69.600 69.200 69.700 ;
        RECT 26.800 67.600 27.600 68.400 ;
        RECT 68.400 68.300 69.200 68.400 ;
        RECT 71.600 68.300 72.400 68.400 ;
        RECT 68.400 67.700 72.400 68.300 ;
        RECT 68.400 67.600 69.200 67.700 ;
        RECT 71.600 67.600 72.400 67.700 ;
        RECT 73.200 68.300 74.000 68.400 ;
        RECT 76.400 68.300 77.200 68.400 ;
        RECT 73.200 67.700 77.200 68.300 ;
        RECT 73.200 67.600 74.000 67.700 ;
        RECT 76.400 67.600 77.200 67.700 ;
        RECT 84.400 68.300 85.200 68.400 ;
        RECT 90.800 68.300 91.600 68.400 ;
        RECT 84.400 67.700 91.600 68.300 ;
        RECT 84.400 67.600 85.200 67.700 ;
        RECT 90.800 67.600 91.600 67.700 ;
        RECT 132.400 68.300 133.200 68.400 ;
        RECT 137.200 68.300 138.000 68.400 ;
        RECT 132.400 67.700 138.000 68.300 ;
        RECT 132.400 67.600 133.200 67.700 ;
        RECT 137.200 67.600 138.000 67.700 ;
        RECT 143.600 68.300 144.400 68.400 ;
        RECT 148.400 68.300 149.200 68.400 ;
        RECT 143.600 67.700 149.200 68.300 ;
        RECT 143.600 67.600 144.400 67.700 ;
        RECT 148.400 67.600 149.200 67.700 ;
        RECT 94.000 66.300 94.800 66.400 ;
        RECT 132.400 66.300 133.200 66.400 ;
        RECT 94.000 65.700 133.200 66.300 ;
        RECT 94.000 65.600 94.800 65.700 ;
        RECT 132.400 65.600 133.200 65.700 ;
        RECT 9.200 64.300 10.000 64.400 ;
        RECT 12.400 64.300 13.200 64.400 ;
        RECT 9.200 63.700 13.200 64.300 ;
        RECT 9.200 63.600 10.000 63.700 ;
        RECT 12.400 63.600 13.200 63.700 ;
        RECT 41.200 64.300 42.000 64.400 ;
        RECT 57.200 64.300 58.000 64.400 ;
        RECT 41.200 63.700 58.000 64.300 ;
        RECT 41.200 63.600 42.000 63.700 ;
        RECT 57.200 63.600 58.000 63.700 ;
        RECT 81.200 64.300 82.000 64.400 ;
        RECT 89.200 64.300 90.000 64.400 ;
        RECT 116.400 64.300 117.200 64.400 ;
        RECT 81.200 63.700 117.200 64.300 ;
        RECT 81.200 63.600 82.000 63.700 ;
        RECT 89.200 63.600 90.000 63.700 ;
        RECT 116.400 63.600 117.200 63.700 ;
        RECT 20.400 62.300 21.200 62.400 ;
        RECT 23.600 62.300 24.400 62.400 ;
        RECT 31.600 62.300 32.400 62.400 ;
        RECT 41.200 62.300 42.000 62.400 ;
        RECT 20.400 61.700 42.000 62.300 ;
        RECT 20.400 61.600 21.200 61.700 ;
        RECT 23.600 61.600 24.400 61.700 ;
        RECT 31.600 61.600 32.400 61.700 ;
        RECT 41.200 61.600 42.000 61.700 ;
        RECT 97.200 59.600 98.000 60.400 ;
        RECT 30.000 58.300 30.800 58.400 ;
        RECT 42.800 58.300 43.600 58.400 ;
        RECT 30.000 57.700 43.600 58.300 ;
        RECT 30.000 57.600 30.800 57.700 ;
        RECT 42.800 57.600 43.600 57.700 ;
        RECT 76.400 58.300 77.200 58.400 ;
        RECT 111.600 58.300 112.400 58.400 ;
        RECT 76.400 57.700 112.400 58.300 ;
        RECT 76.400 57.600 77.200 57.700 ;
        RECT 111.600 57.600 112.400 57.700 ;
        RECT 113.200 57.600 114.000 58.400 ;
        RECT 116.400 58.300 117.200 58.400 ;
        RECT 124.400 58.300 125.200 58.400 ;
        RECT 116.400 57.700 125.200 58.300 ;
        RECT 116.400 57.600 117.200 57.700 ;
        RECT 124.400 57.600 125.200 57.700 ;
        RECT 15.600 56.300 16.400 56.400 ;
        RECT 33.200 56.300 34.000 56.400 ;
        RECT 15.600 55.700 34.000 56.300 ;
        RECT 15.600 55.600 16.400 55.700 ;
        RECT 33.200 55.600 34.000 55.700 ;
        RECT 110.000 56.300 110.800 56.400 ;
        RECT 113.200 56.300 114.000 56.400 ;
        RECT 119.600 56.300 120.400 56.400 ;
        RECT 110.000 55.700 120.400 56.300 ;
        RECT 110.000 55.600 110.800 55.700 ;
        RECT 113.200 55.600 114.000 55.700 ;
        RECT 119.600 55.600 120.400 55.700 ;
        RECT 41.200 54.300 42.000 54.400 ;
        RECT 54.000 54.300 54.800 54.400 ;
        RECT 100.400 54.300 101.200 54.400 ;
        RECT 116.400 54.300 117.200 54.400 ;
        RECT 41.200 53.700 117.200 54.300 ;
        RECT 41.200 53.600 42.000 53.700 ;
        RECT 54.000 53.600 54.800 53.700 ;
        RECT 100.400 53.600 101.200 53.700 ;
        RECT 116.400 53.600 117.200 53.700 ;
        RECT 138.800 54.300 139.600 54.400 ;
        RECT 164.400 54.300 165.200 54.400 ;
        RECT 138.800 53.700 165.200 54.300 ;
        RECT 138.800 53.600 139.600 53.700 ;
        RECT 164.400 53.600 165.200 53.700 ;
        RECT 10.800 52.300 11.600 52.400 ;
        RECT 17.200 52.300 18.000 52.400 ;
        RECT 10.800 51.700 18.000 52.300 ;
        RECT 10.800 51.600 11.600 51.700 ;
        RECT 17.200 51.600 18.000 51.700 ;
        RECT 31.600 52.300 32.400 52.400 ;
        RECT 39.600 52.300 40.400 52.400 ;
        RECT 31.600 51.700 40.400 52.300 ;
        RECT 31.600 51.600 32.400 51.700 ;
        RECT 39.600 51.600 40.400 51.700 ;
        RECT 42.800 52.300 43.600 52.400 ;
        RECT 55.600 52.300 56.400 52.400 ;
        RECT 74.800 52.300 75.600 52.400 ;
        RECT 42.800 51.700 75.600 52.300 ;
        RECT 42.800 51.600 43.600 51.700 ;
        RECT 55.600 51.600 56.400 51.700 ;
        RECT 74.800 51.600 75.600 51.700 ;
        RECT 86.000 52.300 86.800 52.400 ;
        RECT 103.600 52.300 104.400 52.400 ;
        RECT 86.000 51.700 104.400 52.300 ;
        RECT 86.000 51.600 86.800 51.700 ;
        RECT 103.600 51.600 104.400 51.700 ;
        RECT 108.400 52.300 109.200 52.400 ;
        RECT 111.600 52.300 112.400 52.400 ;
        RECT 108.400 51.700 112.400 52.300 ;
        RECT 108.400 51.600 109.200 51.700 ;
        RECT 111.600 51.600 112.400 51.700 ;
        RECT 134.000 52.300 134.800 52.400 ;
        RECT 140.400 52.300 141.200 52.400 ;
        RECT 156.400 52.300 157.200 52.400 ;
        RECT 134.000 51.700 157.200 52.300 ;
        RECT 134.000 51.600 134.800 51.700 ;
        RECT 140.400 51.600 141.200 51.700 ;
        RECT 156.400 51.600 157.200 51.700 ;
        RECT 161.200 51.600 162.000 52.400 ;
        RECT 65.200 50.300 66.000 50.400 ;
        RECT 68.400 50.300 69.200 50.400 ;
        RECT 65.200 49.700 69.200 50.300 ;
        RECT 65.200 49.600 66.000 49.700 ;
        RECT 68.400 49.600 69.200 49.700 ;
        RECT 113.200 50.300 114.000 50.400 ;
        RECT 121.200 50.300 122.000 50.400 ;
        RECT 113.200 49.700 122.000 50.300 ;
        RECT 113.200 49.600 114.000 49.700 ;
        RECT 121.200 49.600 122.000 49.700 ;
        RECT 161.200 50.300 162.000 50.400 ;
        RECT 169.200 50.300 170.000 50.400 ;
        RECT 161.200 49.700 170.000 50.300 ;
        RECT 161.200 49.600 162.000 49.700 ;
        RECT 169.200 49.600 170.000 49.700 ;
        RECT 22.000 48.300 22.800 48.400 ;
        RECT 79.600 48.300 80.400 48.400 ;
        RECT 22.000 47.700 80.400 48.300 ;
        RECT 22.000 47.600 22.800 47.700 ;
        RECT 79.600 47.600 80.400 47.700 ;
        RECT 97.200 48.300 98.000 48.400 ;
        RECT 121.200 48.300 122.000 48.400 ;
        RECT 134.000 48.300 134.800 48.400 ;
        RECT 135.600 48.300 136.400 48.400 ;
        RECT 97.200 47.700 136.400 48.300 ;
        RECT 97.200 47.600 98.000 47.700 ;
        RECT 121.200 47.600 122.000 47.700 ;
        RECT 134.000 47.600 134.800 47.700 ;
        RECT 135.600 47.600 136.400 47.700 ;
        RECT 41.200 46.300 42.000 46.400 ;
        RECT 54.000 46.300 54.800 46.400 ;
        RECT 41.200 45.700 54.800 46.300 ;
        RECT 41.200 45.600 42.000 45.700 ;
        RECT 54.000 45.600 54.800 45.700 ;
        RECT 66.800 46.300 67.600 46.400 ;
        RECT 82.800 46.300 83.600 46.400 ;
        RECT 66.800 45.700 83.600 46.300 ;
        RECT 66.800 45.600 67.600 45.700 ;
        RECT 82.800 45.600 83.600 45.700 ;
        RECT 162.800 46.300 163.600 46.400 ;
        RECT 167.600 46.300 168.400 46.400 ;
        RECT 162.800 45.700 168.400 46.300 ;
        RECT 162.800 45.600 163.600 45.700 ;
        RECT 167.600 45.600 168.400 45.700 ;
        RECT 26.800 44.300 27.600 44.400 ;
        RECT 63.600 44.300 64.400 44.400 ;
        RECT 113.200 44.300 114.000 44.400 ;
        RECT 26.800 43.700 114.000 44.300 ;
        RECT 26.800 43.600 27.600 43.700 ;
        RECT 63.600 43.600 64.400 43.700 ;
        RECT 113.200 43.600 114.000 43.700 ;
        RECT 65.200 42.300 66.000 42.400 ;
        RECT 81.200 42.300 82.000 42.400 ;
        RECT 97.200 42.300 98.000 42.400 ;
        RECT 65.200 41.700 98.000 42.300 ;
        RECT 65.200 41.600 66.000 41.700 ;
        RECT 81.200 41.600 82.000 41.700 ;
        RECT 97.200 41.600 98.000 41.700 ;
        RECT 14.000 38.300 14.800 38.400 ;
        RECT 38.000 38.300 38.800 38.400 ;
        RECT 111.600 38.300 112.400 38.400 ;
        RECT 119.600 38.300 120.400 38.400 ;
        RECT 14.000 37.700 75.500 38.300 ;
        RECT 14.000 37.600 14.800 37.700 ;
        RECT 38.000 37.600 38.800 37.700 ;
        RECT 74.900 36.400 75.500 37.700 ;
        RECT 111.600 37.700 120.400 38.300 ;
        RECT 111.600 37.600 112.400 37.700 ;
        RECT 119.600 37.600 120.400 37.700 ;
        RECT 31.600 36.300 32.400 36.400 ;
        RECT 41.200 36.300 42.000 36.400 ;
        RECT 31.600 35.700 42.000 36.300 ;
        RECT 31.600 35.600 32.400 35.700 ;
        RECT 41.200 35.600 42.000 35.700 ;
        RECT 74.800 36.300 75.600 36.400 ;
        RECT 92.400 36.300 93.200 36.400 ;
        RECT 74.800 35.700 93.200 36.300 ;
        RECT 74.800 35.600 75.600 35.700 ;
        RECT 92.400 35.600 93.200 35.700 ;
        RECT 34.800 34.300 35.600 34.400 ;
        RECT 46.000 34.300 46.800 34.400 ;
        RECT 105.200 34.300 106.000 34.400 ;
        RECT 34.800 33.700 106.000 34.300 ;
        RECT 34.800 33.600 35.600 33.700 ;
        RECT 46.000 33.600 46.800 33.700 ;
        RECT 105.200 33.600 106.000 33.700 ;
        RECT 9.200 32.300 10.000 32.400 ;
        RECT 25.200 32.300 26.000 32.400 ;
        RECT 9.200 31.700 26.000 32.300 ;
        RECT 9.200 31.600 10.000 31.700 ;
        RECT 25.200 31.600 26.000 31.700 ;
        RECT 42.800 32.300 43.600 32.400 ;
        RECT 76.400 32.300 77.200 32.400 ;
        RECT 42.800 31.700 77.200 32.300 ;
        RECT 42.800 31.600 43.600 31.700 ;
        RECT 76.400 31.600 77.200 31.700 ;
        RECT 102.000 32.300 102.800 32.400 ;
        RECT 106.800 32.300 107.600 32.400 ;
        RECT 102.000 31.700 107.600 32.300 ;
        RECT 102.000 31.600 102.800 31.700 ;
        RECT 106.800 31.600 107.600 31.700 ;
        RECT 111.600 32.300 112.400 32.400 ;
        RECT 113.200 32.300 114.000 32.400 ;
        RECT 111.600 31.700 114.000 32.300 ;
        RECT 111.600 31.600 112.400 31.700 ;
        RECT 113.200 31.600 114.000 31.700 ;
        RECT 7.600 30.300 8.400 30.400 ;
        RECT 15.600 30.300 16.400 30.400 ;
        RECT 7.600 29.700 16.400 30.300 ;
        RECT 7.600 29.600 8.400 29.700 ;
        RECT 15.600 29.600 16.400 29.700 ;
        RECT 39.600 30.300 40.400 30.400 ;
        RECT 78.000 30.300 78.800 30.400 ;
        RECT 39.600 29.700 78.800 30.300 ;
        RECT 39.600 29.600 40.400 29.700 ;
        RECT 78.000 29.600 78.800 29.700 ;
        RECT 79.600 30.300 80.400 30.400 ;
        RECT 90.800 30.300 91.600 30.400 ;
        RECT 103.600 30.300 104.400 30.400 ;
        RECT 79.600 29.700 104.400 30.300 ;
        RECT 79.600 29.600 80.400 29.700 ;
        RECT 90.800 29.600 91.600 29.700 ;
        RECT 103.600 29.600 104.400 29.700 ;
        RECT 105.200 30.300 106.000 30.400 ;
        RECT 113.200 30.300 114.000 30.400 ;
        RECT 105.200 29.700 114.000 30.300 ;
        RECT 105.200 29.600 106.000 29.700 ;
        RECT 113.200 29.600 114.000 29.700 ;
        RECT 118.000 30.300 118.800 30.400 ;
        RECT 129.200 30.300 130.000 30.400 ;
        RECT 118.000 29.700 130.000 30.300 ;
        RECT 118.000 29.600 118.800 29.700 ;
        RECT 129.200 29.600 130.000 29.700 ;
        RECT 140.400 30.300 141.200 30.400 ;
        RECT 161.200 30.300 162.000 30.400 ;
        RECT 162.800 30.300 163.600 30.400 ;
        RECT 140.400 29.700 163.600 30.300 ;
        RECT 140.400 29.600 141.200 29.700 ;
        RECT 161.200 29.600 162.000 29.700 ;
        RECT 162.800 29.600 163.600 29.700 ;
        RECT 17.200 28.300 18.000 28.400 ;
        RECT 22.000 28.300 22.800 28.400 ;
        RECT 38.000 28.300 38.800 28.400 ;
        RECT 17.200 27.700 38.800 28.300 ;
        RECT 17.200 27.600 18.000 27.700 ;
        RECT 22.000 27.600 22.800 27.700 ;
        RECT 38.000 27.600 38.800 27.700 ;
        RECT 76.400 28.300 77.200 28.400 ;
        RECT 81.200 28.300 82.000 28.400 ;
        RECT 76.400 27.700 82.000 28.300 ;
        RECT 76.400 27.600 77.200 27.700 ;
        RECT 81.200 27.600 82.000 27.700 ;
        RECT 135.600 28.300 136.400 28.400 ;
        RECT 146.800 28.300 147.600 28.400 ;
        RECT 135.600 27.700 147.600 28.300 ;
        RECT 135.600 27.600 136.400 27.700 ;
        RECT 146.800 27.600 147.600 27.700 ;
        RECT 20.400 26.300 21.200 26.400 ;
        RECT 26.800 26.300 27.600 26.400 ;
        RECT 20.400 25.700 27.600 26.300 ;
        RECT 20.400 25.600 21.200 25.700 ;
        RECT 26.800 25.600 27.600 25.700 ;
        RECT 97.200 24.300 98.000 24.400 ;
        RECT 135.600 24.300 136.400 24.400 ;
        RECT 140.400 24.300 141.200 24.400 ;
        RECT 158.000 24.300 158.800 24.400 ;
        RECT 159.600 24.300 160.400 24.400 ;
        RECT 97.200 23.700 160.400 24.300 ;
        RECT 97.200 23.600 98.000 23.700 ;
        RECT 135.600 23.600 136.400 23.700 ;
        RECT 140.400 23.600 141.200 23.700 ;
        RECT 158.000 23.600 158.800 23.700 ;
        RECT 159.600 23.600 160.400 23.700 ;
        RECT 161.200 24.300 162.000 24.400 ;
        RECT 170.800 24.300 171.600 24.400 ;
        RECT 161.200 23.700 171.600 24.300 ;
        RECT 161.200 23.600 162.000 23.700 ;
        RECT 170.800 23.600 171.600 23.700 ;
        RECT 169.200 22.300 170.000 22.400 ;
        RECT 177.200 22.300 178.000 22.400 ;
        RECT 169.200 21.700 178.000 22.300 ;
        RECT 169.200 21.600 170.000 21.700 ;
        RECT 177.200 21.600 178.000 21.700 ;
        RECT 10.800 18.300 11.600 18.400 ;
        RECT 26.800 18.300 27.600 18.400 ;
        RECT 44.400 18.300 45.200 18.400 ;
        RECT 68.400 18.300 69.200 18.400 ;
        RECT 89.200 18.300 90.000 18.400 ;
        RECT 97.200 18.300 98.000 18.400 ;
        RECT 10.800 17.700 98.000 18.300 ;
        RECT 10.800 17.600 11.600 17.700 ;
        RECT 26.800 17.600 27.600 17.700 ;
        RECT 44.400 17.600 45.200 17.700 ;
        RECT 68.400 17.600 69.200 17.700 ;
        RECT 89.200 17.600 90.000 17.700 ;
        RECT 97.200 17.600 98.000 17.700 ;
        RECT 106.800 18.300 107.600 18.400 ;
        RECT 111.600 18.300 112.400 18.400 ;
        RECT 114.800 18.300 115.600 18.400 ;
        RECT 106.800 17.700 110.700 18.300 ;
        RECT 106.800 17.600 107.600 17.700 ;
        RECT 71.600 16.300 72.400 16.400 ;
        RECT 76.400 16.300 77.200 16.400 ;
        RECT 97.200 16.300 98.000 16.400 ;
        RECT 71.600 15.700 98.000 16.300 ;
        RECT 110.100 16.300 110.700 17.700 ;
        RECT 111.600 17.700 115.600 18.300 ;
        RECT 111.600 17.600 112.400 17.700 ;
        RECT 114.800 17.600 115.600 17.700 ;
        RECT 159.600 16.300 160.400 16.400 ;
        RECT 110.100 15.700 160.400 16.300 ;
        RECT 71.600 15.600 72.400 15.700 ;
        RECT 76.400 15.600 77.200 15.700 ;
        RECT 97.200 15.600 98.000 15.700 ;
        RECT 159.600 15.600 160.400 15.700 ;
        RECT 14.000 14.300 14.800 14.400 ;
        RECT 22.000 14.300 22.800 14.400 ;
        RECT 14.000 13.700 22.800 14.300 ;
        RECT 14.000 13.600 14.800 13.700 ;
        RECT 22.000 13.600 22.800 13.700 ;
        RECT 42.800 14.300 43.600 14.400 ;
        RECT 46.000 14.300 46.800 14.400 ;
        RECT 78.000 14.300 78.800 14.400 ;
        RECT 42.800 13.700 46.800 14.300 ;
        RECT 42.800 13.600 43.600 13.700 ;
        RECT 46.000 13.600 46.800 13.700 ;
        RECT 47.700 13.700 78.800 14.300 ;
        RECT 14.000 11.600 14.800 12.400 ;
        RECT 15.600 12.300 16.400 12.400 ;
        RECT 26.800 12.300 27.600 12.400 ;
        RECT 44.400 12.300 45.200 12.400 ;
        RECT 47.700 12.300 48.300 13.700 ;
        RECT 78.000 13.600 78.800 13.700 ;
        RECT 129.200 14.300 130.000 14.400 ;
        RECT 135.600 14.300 136.400 14.400 ;
        RECT 129.200 13.700 136.400 14.300 ;
        RECT 129.200 13.600 130.000 13.700 ;
        RECT 135.600 13.600 136.400 13.700 ;
        RECT 172.400 14.300 173.200 14.400 ;
        RECT 175.600 14.300 176.400 14.400 ;
        RECT 172.400 13.700 176.400 14.300 ;
        RECT 172.400 13.600 173.200 13.700 ;
        RECT 175.600 13.600 176.400 13.700 ;
        RECT 15.600 11.700 48.300 12.300 ;
        RECT 63.600 12.300 64.400 12.400 ;
        RECT 70.000 12.300 70.800 12.400 ;
        RECT 73.200 12.300 74.000 12.400 ;
        RECT 63.600 11.700 74.000 12.300 ;
        RECT 15.600 11.600 16.400 11.700 ;
        RECT 26.800 11.600 27.600 11.700 ;
        RECT 44.400 11.600 45.200 11.700 ;
        RECT 63.600 11.600 64.400 11.700 ;
        RECT 70.000 11.600 70.800 11.700 ;
        RECT 73.200 11.600 74.000 11.700 ;
        RECT 81.200 12.300 82.000 12.400 ;
        RECT 84.400 12.300 85.200 12.400 ;
        RECT 81.200 11.700 85.200 12.300 ;
        RECT 81.200 11.600 82.000 11.700 ;
        RECT 84.400 11.600 85.200 11.700 ;
        RECT 132.400 12.300 133.200 12.400 ;
        RECT 140.400 12.300 141.200 12.400 ;
        RECT 132.400 11.700 141.200 12.300 ;
        RECT 132.400 11.600 133.200 11.700 ;
        RECT 140.400 11.600 141.200 11.700 ;
        RECT 142.000 12.300 142.800 12.400 ;
        RECT 145.200 12.300 146.000 12.400 ;
        RECT 142.000 11.700 146.000 12.300 ;
        RECT 142.000 11.600 142.800 11.700 ;
        RECT 145.200 11.600 146.000 11.700 ;
        RECT 154.800 12.300 155.600 12.400 ;
        RECT 162.800 12.300 163.600 12.400 ;
        RECT 154.800 11.700 163.600 12.300 ;
        RECT 154.800 11.600 155.600 11.700 ;
        RECT 162.800 11.600 163.600 11.700 ;
      LAYER metal4 ;
        RECT 4.200 71.400 5.400 96.600 ;
        RECT 26.600 43.400 27.800 68.600 ;
        RECT 13.800 11.400 15.000 38.600 ;
        RECT 77.800 29.400 79.000 72.600 ;
        RECT 81.000 11.400 82.200 42.600 ;
        RECT 97.000 17.400 98.200 100.600 ;
        RECT 113.000 31.400 114.200 58.600 ;
        RECT 161.000 23.400 162.200 52.600 ;
  END
END sigmoid_approx
END LIBRARY

