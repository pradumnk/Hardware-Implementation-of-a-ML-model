magic
tech scmos
magscale 1 2
timestamp 1646624542
<< checkpaint >>
rect -544 -400 556 936
<< metal1 >>
rect -442 870 -374 872
rect -442 862 -439 870
rect -421 862 -374 870
rect -442 860 -374 862
rect -484 670 -374 672
rect -484 662 -481 670
rect -463 662 -374 670
rect -484 660 -374 662
rect -442 630 -390 632
rect -442 622 -439 630
rect -421 622 -390 630
rect -442 620 -390 622
rect -484 430 -392 432
rect -484 422 -481 430
rect -463 422 -392 430
rect -484 420 -392 422
rect -442 402 -380 404
rect -442 394 -439 402
rect -421 394 -380 402
rect -442 392 -380 394
rect -484 202 -376 204
rect -484 194 -481 202
rect -463 194 -376 202
rect -484 192 -376 194
rect -442 152 -374 154
rect -442 144 -439 152
rect -421 144 -374 152
rect -442 142 -374 144
rect -484 -48 -374 -46
rect -484 -56 -481 -48
rect -463 -56 -374 -48
rect -484 -58 -374 -56
rect -442 -96 -348 -94
rect -442 -104 -439 -96
rect -421 -104 -348 -96
rect -442 -106 -348 -104
rect -484 -296 -348 -294
rect -484 -304 -481 -296
rect -463 -304 -348 -296
rect -484 -306 -348 -304
<< m2contact >>
rect -439 862 -421 870
rect -481 662 -463 670
rect -439 622 -421 630
rect -481 422 -463 430
rect -439 394 -421 402
rect -481 194 -463 202
rect -439 144 -421 152
rect -481 -56 -463 -48
rect -439 -104 -421 -96
rect -481 -304 -463 -296
<< metal2 >>
rect -442 870 -418 872
rect -442 862 -439 870
rect -421 862 -418 870
rect -484 670 -460 672
rect -484 662 -481 670
rect -463 662 -460 670
rect -484 430 -460 662
rect -484 422 -481 430
rect -463 422 -460 430
rect -484 202 -460 422
rect -484 194 -481 202
rect -463 194 -460 202
rect -484 -48 -460 194
rect -484 -56 -481 -48
rect -463 -56 -460 -48
rect -484 -296 -460 -56
rect -484 -304 -481 -296
rect -463 -304 -460 -296
rect -484 -340 -460 -304
rect -442 630 -418 862
rect -442 622 -439 630
rect -421 622 -418 630
rect -442 402 -418 622
rect -442 394 -439 402
rect -421 394 -418 402
rect -442 152 -418 394
rect -442 144 -439 152
rect -421 144 -418 152
rect -442 -96 -418 144
rect -442 -104 -439 -96
rect -421 -104 -418 -96
rect -442 -340 -418 -104
use CLKBUF3  CLKBUF3_0
timestamp 1646624542
transform 1 0 0 0 1 -300
box -16 -6 288 210
use CLKBUF2  CLKBUF2_0
timestamp 1646624542
transform 1 0 -208 0 1 -300
box -16 -6 224 210
use CLKBUF1  CLKBUF1_0
timestamp 1646624542
transform 1 0 -352 0 1 -300
box -16 -6 160 210
use DFFSR  DFFSR_0
timestamp 1646624542
transform 1 0 -148 0 1 -52
box -16 -6 368 210
use LATCH  LATCH_0
timestamp 1646624542
transform 1 0 -260 0 1 -52
box -16 -6 128 210
use XNOR2X1  XNOR2X1_0
timestamp 1646624542
transform 1 0 -372 0 1 -52
box -16 -6 128 210
use MUX2X1  MUX2X1_0
timestamp 1646624542
transform 1 0 390 0 1 198
box -10 -6 106 210
use XOR2X1  XOR2X1_0
timestamp 1646624542
transform 1 0 278 0 1 198
box -16 -6 128 210
use TBUFX2  TBUFX2_0
timestamp 1646624542
transform 1 0 162 0 1 198
box -10 -6 120 210
use TBUFX1  TBUFX1_0
timestamp 1646624542
transform 1 0 82 0 1 198
box -10 -6 84 210
use OR2X2  OR2X2_0
timestamp 1646624542
transform 1 0 10 0 1 198
box -14 -6 70 210
use OR2X1  OR2X1_0
timestamp 1646624542
transform 1 0 -58 0 1 198
box -16 -6 80 210
use OAI22X1  OAI22X1_0
timestamp 1646624542
transform 1 0 -146 0 1 198
box -16 -6 92 210
use OAI21X1  OAI21X1_0
timestamp 1646624542
transform 1 0 -218 0 1 198
box -16 -6 68 210
use NOR2X1  NOR2X1_0
timestamp 1646624542
transform 1 0 -270 0 1 198
box -16 -6 64 210
use NAND3X1  NAND3X1_0
timestamp 1646624542
transform 1 0 -340 0 1 198
box -16 -6 80 210
use NAND2X1  NAND2X1_0
timestamp 1646624542
transform 1 0 -388 0 1 198
box -16 -6 64 210
use INVX8  INVX8_0
timestamp 1646624542
transform 1 0 322 0 1 426
box -18 -6 90 210
use INVX4  INVX4_0
timestamp 1646624542
transform 1 0 274 0 1 426
box -18 -6 56 210
use INVX2  INVX2_0
timestamp 1646624542
transform 1 0 242 0 1 426
box -18 -6 52 210
use INVX1  INVX1_0
timestamp 1646624542
transform 1 0 210 0 1 426
box -18 -6 52 210
use HAX1  HAX1_0
timestamp 1646624542
transform 1 0 44 0 1 426
box -10 -6 168 210
use FAX1  FAX1_0
timestamp 1646624542
transform 1 0 -202 0 1 426
box -10 -6 252 210
use DFFPOSX1  DFFPOSX1_0
timestamp 1646624542
transform 1 0 -400 0 1 426
box -16 -6 208 210
use NOR3X1  NOR3X1_0
timestamp 1646624542
transform 1 0 228 0 1 666
box -14 -6 136 210
use DFFNEGX1  DFFNEGX1_0
timestamp 1646624542
transform 1 0 32 0 1 666
box -16 -6 208 210
use BUFX4  BUFX4_0
timestamp 1646624542
transform 1 0 -38 0 1 666
box -18 -6 74 210
use BUFX2  BUFX2_0
timestamp 1646624542
transform 1 0 -86 0 1 666
box -10 -6 56 210
use AOI22X1  AOI22X1_0
timestamp 1646624542
transform 1 0 -168 0 1 666
box -16 -6 92 210
use AOI21X1  AOI21X1_0
timestamp 1646624542
transform 1 0 -232 0 1 666
box -14 -6 78 210
use AND2X2  AND2X2_0
timestamp 1646624542
transform 1 0 -298 0 1 666
box -16 -6 80 210
use AND2X1  AND2X1_0
timestamp 1646624542
transform 1 0 -362 0 1 666
box -16 -6 80 210
use FILL  FILL_0
timestamp 1646624542
transform 1 0 -378 0 1 666
box -16 -6 32 210
<< end >>
