magic
tech scmos
magscale 1 2
timestamp 1646624542
<< checkpaint >>
rect -70 -66 180 270
<< nwell >>
rect -10 96 120 210
<< ntransistor >>
rect 14 12 18 52
rect 46 12 50 52
rect 62 12 66 52
rect 78 12 82 52
rect 94 12 98 52
<< ptransistor >>
rect 14 108 18 188
rect 46 108 50 188
rect 62 108 66 188
rect 78 108 82 188
rect 94 108 98 188
<< ndiffusion >>
rect 4 51 14 52
rect 12 13 14 51
rect 4 12 14 13
rect 18 51 28 52
rect 18 13 20 51
rect 18 12 28 13
rect 36 51 46 52
rect 44 13 46 51
rect 36 12 46 13
rect 50 24 52 52
rect 60 24 62 52
rect 50 12 62 24
rect 66 51 78 52
rect 66 13 68 51
rect 76 13 78 51
rect 66 12 78 13
rect 82 43 94 52
rect 82 15 84 43
rect 92 15 94 43
rect 82 12 94 15
rect 98 43 108 52
rect 98 15 100 43
rect 98 12 108 15
<< pdiffusion >>
rect 4 187 14 188
rect 12 109 14 187
rect 4 108 14 109
rect 18 187 28 188
rect 18 109 20 187
rect 18 108 28 109
rect 36 187 46 188
rect 44 109 46 187
rect 36 108 46 109
rect 50 176 62 188
rect 50 108 52 176
rect 60 108 62 176
rect 66 187 78 188
rect 66 109 68 187
rect 76 109 78 187
rect 66 108 78 109
rect 82 184 94 188
rect 82 126 84 184
rect 92 126 94 184
rect 82 108 94 126
rect 98 187 108 188
rect 98 109 100 187
rect 98 108 108 109
<< ndcontact >>
rect 4 13 12 51
rect 20 13 28 51
rect 36 13 44 51
rect 52 24 60 52
rect 68 13 76 51
rect 84 15 92 43
rect 100 15 108 43
<< pdcontact >>
rect 4 109 12 187
rect 20 109 28 187
rect 36 109 44 187
rect 52 108 60 176
rect 68 109 76 187
rect 84 126 92 184
rect 100 109 108 187
<< psubstratepcontact >>
rect -4 -4 4 4
rect 28 -4 36 4
rect 60 -4 68 4
rect 92 -4 100 4
<< nsubstratencontact >>
rect -4 196 4 204
rect 28 196 36 204
rect 60 196 68 204
rect 92 196 100 204
<< polysilicon >>
rect 14 188 18 192
rect 46 188 50 192
rect 62 188 66 192
rect 78 188 82 192
rect 94 188 98 192
rect 14 102 18 108
rect 46 106 50 108
rect 62 106 66 108
rect 12 98 18 102
rect 24 102 66 106
rect 78 106 82 108
rect 94 106 98 108
rect 78 102 98 106
rect 24 90 28 102
rect 94 74 98 102
rect 14 58 18 66
rect 94 58 98 66
rect 14 54 66 58
rect 14 52 18 54
rect 46 52 50 54
rect 62 52 66 54
rect 78 54 98 58
rect 78 52 82 54
rect 94 52 98 54
rect 14 8 18 12
rect 46 8 50 12
rect 62 8 66 12
rect 78 8 82 12
rect 94 8 98 12
<< polycontact >>
rect 4 94 12 102
rect 20 82 28 90
rect 90 66 98 74
rect 6 58 14 66
<< metal1 >>
rect -4 204 116 206
rect 4 196 28 204
rect 36 196 60 204
rect 68 196 92 204
rect 100 196 116 204
rect -4 194 116 196
rect 4 187 12 194
rect 4 108 12 109
rect 20 187 28 188
rect 20 108 28 109
rect 36 187 76 188
rect 44 182 68 187
rect 36 108 44 109
rect 84 184 92 194
rect 84 122 92 126
rect 100 187 108 188
rect 76 109 100 116
rect 68 108 108 109
rect 4 86 12 94
rect 20 90 26 108
rect 52 94 58 108
rect 4 66 10 86
rect 52 86 60 94
rect 4 58 6 66
rect 20 52 26 82
rect 52 52 58 86
rect 98 66 108 74
rect 68 52 108 58
rect 4 51 12 52
rect 4 6 12 13
rect 20 51 28 52
rect 20 12 28 13
rect 36 51 44 52
rect 68 51 76 52
rect 44 13 68 18
rect 102 46 108 52
rect 36 12 76 13
rect 84 43 92 46
rect 84 6 92 15
rect 100 43 108 46
rect 100 12 108 15
rect -4 4 116 6
rect 4 -4 28 4
rect 36 -4 60 4
rect 68 -4 92 4
rect 100 -4 116 4
rect -4 -6 116 -4
<< m1p >>
rect 4 86 12 94
rect 52 86 60 94
rect 100 66 108 74
<< labels >>
rlabel metal1 8 200 8 200 4 vdd
rlabel metal1 8 0 8 0 4 gnd
rlabel metal1 104 70 104 70 4 A
rlabel metal1 8 90 8 90 4 EN
rlabel metal1 56 90 56 90 4 Y
<< end >>
